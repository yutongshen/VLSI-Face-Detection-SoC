../include/CtrlSignal.svh