PLIC/Target.sv