AHB/MuxM2S.sv