../include/Interrupt_def.svh