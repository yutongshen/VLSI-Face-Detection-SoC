../include/FunctCode.svh