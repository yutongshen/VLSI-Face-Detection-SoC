../include/ForwardCtrl.svh