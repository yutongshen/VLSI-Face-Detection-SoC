../include/OPCode.svh