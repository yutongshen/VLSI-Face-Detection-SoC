# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SRAM_small
#       Words            : 512
#       Bits             : 8
#       Byte-Write       : 4
#       Aspect Ratio     : 1
#       Output Loading   : 0.01  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2019/01/14 16:00:55
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SRAM_small
CLASS BLOCK ;
FOREIGN SRAM_small 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 553.040 BY 294.000 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 551.920 282.580 553.040 285.820 ;
  LAYER ME3 ;
  RECT 551.920 282.580 553.040 285.820 ;
  LAYER ME2 ;
  RECT 551.920 282.580 553.040 285.820 ;
  LAYER ME1 ;
  RECT 551.920 282.580 553.040 285.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 274.740 553.040 277.980 ;
  LAYER ME3 ;
  RECT 551.920 274.740 553.040 277.980 ;
  LAYER ME2 ;
  RECT 551.920 274.740 553.040 277.980 ;
  LAYER ME1 ;
  RECT 551.920 274.740 553.040 277.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 266.900 553.040 270.140 ;
  LAYER ME3 ;
  RECT 551.920 266.900 553.040 270.140 ;
  LAYER ME2 ;
  RECT 551.920 266.900 553.040 270.140 ;
  LAYER ME1 ;
  RECT 551.920 266.900 553.040 270.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 259.060 553.040 262.300 ;
  LAYER ME3 ;
  RECT 551.920 259.060 553.040 262.300 ;
  LAYER ME2 ;
  RECT 551.920 259.060 553.040 262.300 ;
  LAYER ME1 ;
  RECT 551.920 259.060 553.040 262.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 251.220 553.040 254.460 ;
  LAYER ME3 ;
  RECT 551.920 251.220 553.040 254.460 ;
  LAYER ME2 ;
  RECT 551.920 251.220 553.040 254.460 ;
  LAYER ME1 ;
  RECT 551.920 251.220 553.040 254.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 243.380 553.040 246.620 ;
  LAYER ME3 ;
  RECT 551.920 243.380 553.040 246.620 ;
  LAYER ME2 ;
  RECT 551.920 243.380 553.040 246.620 ;
  LAYER ME1 ;
  RECT 551.920 243.380 553.040 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 204.180 553.040 207.420 ;
  LAYER ME3 ;
  RECT 551.920 204.180 553.040 207.420 ;
  LAYER ME2 ;
  RECT 551.920 204.180 553.040 207.420 ;
  LAYER ME1 ;
  RECT 551.920 204.180 553.040 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 196.340 553.040 199.580 ;
  LAYER ME3 ;
  RECT 551.920 196.340 553.040 199.580 ;
  LAYER ME2 ;
  RECT 551.920 196.340 553.040 199.580 ;
  LAYER ME1 ;
  RECT 551.920 196.340 553.040 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 188.500 553.040 191.740 ;
  LAYER ME3 ;
  RECT 551.920 188.500 553.040 191.740 ;
  LAYER ME2 ;
  RECT 551.920 188.500 553.040 191.740 ;
  LAYER ME1 ;
  RECT 551.920 188.500 553.040 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 180.660 553.040 183.900 ;
  LAYER ME3 ;
  RECT 551.920 180.660 553.040 183.900 ;
  LAYER ME2 ;
  RECT 551.920 180.660 553.040 183.900 ;
  LAYER ME1 ;
  RECT 551.920 180.660 553.040 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 172.820 553.040 176.060 ;
  LAYER ME3 ;
  RECT 551.920 172.820 553.040 176.060 ;
  LAYER ME2 ;
  RECT 551.920 172.820 553.040 176.060 ;
  LAYER ME1 ;
  RECT 551.920 172.820 553.040 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 164.980 553.040 168.220 ;
  LAYER ME3 ;
  RECT 551.920 164.980 553.040 168.220 ;
  LAYER ME2 ;
  RECT 551.920 164.980 553.040 168.220 ;
  LAYER ME1 ;
  RECT 551.920 164.980 553.040 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 125.780 553.040 129.020 ;
  LAYER ME3 ;
  RECT 551.920 125.780 553.040 129.020 ;
  LAYER ME2 ;
  RECT 551.920 125.780 553.040 129.020 ;
  LAYER ME1 ;
  RECT 551.920 125.780 553.040 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 117.940 553.040 121.180 ;
  LAYER ME3 ;
  RECT 551.920 117.940 553.040 121.180 ;
  LAYER ME2 ;
  RECT 551.920 117.940 553.040 121.180 ;
  LAYER ME1 ;
  RECT 551.920 117.940 553.040 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 110.100 553.040 113.340 ;
  LAYER ME3 ;
  RECT 551.920 110.100 553.040 113.340 ;
  LAYER ME2 ;
  RECT 551.920 110.100 553.040 113.340 ;
  LAYER ME1 ;
  RECT 551.920 110.100 553.040 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 102.260 553.040 105.500 ;
  LAYER ME3 ;
  RECT 551.920 102.260 553.040 105.500 ;
  LAYER ME2 ;
  RECT 551.920 102.260 553.040 105.500 ;
  LAYER ME1 ;
  RECT 551.920 102.260 553.040 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 94.420 553.040 97.660 ;
  LAYER ME3 ;
  RECT 551.920 94.420 553.040 97.660 ;
  LAYER ME2 ;
  RECT 551.920 94.420 553.040 97.660 ;
  LAYER ME1 ;
  RECT 551.920 94.420 553.040 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 86.580 553.040 89.820 ;
  LAYER ME3 ;
  RECT 551.920 86.580 553.040 89.820 ;
  LAYER ME2 ;
  RECT 551.920 86.580 553.040 89.820 ;
  LAYER ME1 ;
  RECT 551.920 86.580 553.040 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 47.380 553.040 50.620 ;
  LAYER ME3 ;
  RECT 551.920 47.380 553.040 50.620 ;
  LAYER ME2 ;
  RECT 551.920 47.380 553.040 50.620 ;
  LAYER ME1 ;
  RECT 551.920 47.380 553.040 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 39.540 553.040 42.780 ;
  LAYER ME3 ;
  RECT 551.920 39.540 553.040 42.780 ;
  LAYER ME2 ;
  RECT 551.920 39.540 553.040 42.780 ;
  LAYER ME1 ;
  RECT 551.920 39.540 553.040 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 31.700 553.040 34.940 ;
  LAYER ME3 ;
  RECT 551.920 31.700 553.040 34.940 ;
  LAYER ME2 ;
  RECT 551.920 31.700 553.040 34.940 ;
  LAYER ME1 ;
  RECT 551.920 31.700 553.040 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 23.860 553.040 27.100 ;
  LAYER ME3 ;
  RECT 551.920 23.860 553.040 27.100 ;
  LAYER ME2 ;
  RECT 551.920 23.860 553.040 27.100 ;
  LAYER ME1 ;
  RECT 551.920 23.860 553.040 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 16.020 553.040 19.260 ;
  LAYER ME3 ;
  RECT 551.920 16.020 553.040 19.260 ;
  LAYER ME2 ;
  RECT 551.920 16.020 553.040 19.260 ;
  LAYER ME1 ;
  RECT 551.920 16.020 553.040 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 8.180 553.040 11.420 ;
  LAYER ME3 ;
  RECT 551.920 8.180 553.040 11.420 ;
  LAYER ME2 ;
  RECT 551.920 8.180 553.040 11.420 ;
  LAYER ME1 ;
  RECT 551.920 8.180 553.040 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.320 292.880 540.860 294.000 ;
  LAYER ME3 ;
  RECT 537.320 292.880 540.860 294.000 ;
  LAYER ME2 ;
  RECT 537.320 292.880 540.860 294.000 ;
  LAYER ME1 ;
  RECT 537.320 292.880 540.860 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.640 292.880 532.180 294.000 ;
  LAYER ME3 ;
  RECT 528.640 292.880 532.180 294.000 ;
  LAYER ME2 ;
  RECT 528.640 292.880 532.180 294.000 ;
  LAYER ME1 ;
  RECT 528.640 292.880 532.180 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.240 292.880 488.780 294.000 ;
  LAYER ME3 ;
  RECT 485.240 292.880 488.780 294.000 ;
  LAYER ME2 ;
  RECT 485.240 292.880 488.780 294.000 ;
  LAYER ME1 ;
  RECT 485.240 292.880 488.780 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.560 292.880 480.100 294.000 ;
  LAYER ME3 ;
  RECT 476.560 292.880 480.100 294.000 ;
  LAYER ME2 ;
  RECT 476.560 292.880 480.100 294.000 ;
  LAYER ME1 ;
  RECT 476.560 292.880 480.100 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.880 292.880 471.420 294.000 ;
  LAYER ME3 ;
  RECT 467.880 292.880 471.420 294.000 ;
  LAYER ME2 ;
  RECT 467.880 292.880 471.420 294.000 ;
  LAYER ME1 ;
  RECT 467.880 292.880 471.420 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.200 292.880 462.740 294.000 ;
  LAYER ME3 ;
  RECT 459.200 292.880 462.740 294.000 ;
  LAYER ME2 ;
  RECT 459.200 292.880 462.740 294.000 ;
  LAYER ME1 ;
  RECT 459.200 292.880 462.740 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.520 292.880 454.060 294.000 ;
  LAYER ME3 ;
  RECT 450.520 292.880 454.060 294.000 ;
  LAYER ME2 ;
  RECT 450.520 292.880 454.060 294.000 ;
  LAYER ME1 ;
  RECT 450.520 292.880 454.060 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.840 292.880 445.380 294.000 ;
  LAYER ME3 ;
  RECT 441.840 292.880 445.380 294.000 ;
  LAYER ME2 ;
  RECT 441.840 292.880 445.380 294.000 ;
  LAYER ME1 ;
  RECT 441.840 292.880 445.380 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.440 292.880 401.980 294.000 ;
  LAYER ME3 ;
  RECT 398.440 292.880 401.980 294.000 ;
  LAYER ME2 ;
  RECT 398.440 292.880 401.980 294.000 ;
  LAYER ME1 ;
  RECT 398.440 292.880 401.980 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.760 292.880 393.300 294.000 ;
  LAYER ME3 ;
  RECT 389.760 292.880 393.300 294.000 ;
  LAYER ME2 ;
  RECT 389.760 292.880 393.300 294.000 ;
  LAYER ME1 ;
  RECT 389.760 292.880 393.300 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.080 292.880 384.620 294.000 ;
  LAYER ME3 ;
  RECT 381.080 292.880 384.620 294.000 ;
  LAYER ME2 ;
  RECT 381.080 292.880 384.620 294.000 ;
  LAYER ME1 ;
  RECT 381.080 292.880 384.620 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.400 292.880 375.940 294.000 ;
  LAYER ME3 ;
  RECT 372.400 292.880 375.940 294.000 ;
  LAYER ME2 ;
  RECT 372.400 292.880 375.940 294.000 ;
  LAYER ME1 ;
  RECT 372.400 292.880 375.940 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 292.880 367.260 294.000 ;
  LAYER ME3 ;
  RECT 363.720 292.880 367.260 294.000 ;
  LAYER ME2 ;
  RECT 363.720 292.880 367.260 294.000 ;
  LAYER ME1 ;
  RECT 363.720 292.880 367.260 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.040 292.880 358.580 294.000 ;
  LAYER ME3 ;
  RECT 355.040 292.880 358.580 294.000 ;
  LAYER ME2 ;
  RECT 355.040 292.880 358.580 294.000 ;
  LAYER ME1 ;
  RECT 355.040 292.880 358.580 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER ME3 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER ME2 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER ME1 ;
  RECT 311.640 292.880 315.180 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER ME3 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER ME2 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER ME1 ;
  RECT 302.960 292.880 306.500 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER ME3 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER ME2 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER ME1 ;
  RECT 294.280 292.880 297.820 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER ME3 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER ME2 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER ME1 ;
  RECT 285.600 292.880 289.140 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER ME3 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER ME2 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER ME1 ;
  RECT 276.920 292.880 280.460 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER ME3 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER ME2 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER ME1 ;
  RECT 268.240 292.880 271.780 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER ME3 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER ME2 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER ME1 ;
  RECT 224.840 292.880 228.380 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER ME3 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER ME2 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER ME1 ;
  RECT 216.160 292.880 219.700 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER ME3 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER ME2 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER ME1 ;
  RECT 207.480 292.880 211.020 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER ME3 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER ME2 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER ME1 ;
  RECT 198.800 292.880 202.340 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER ME3 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER ME2 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER ME1 ;
  RECT 190.120 292.880 193.660 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER ME3 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER ME2 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER ME1 ;
  RECT 181.440 292.880 184.980 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER ME3 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER ME2 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER ME1 ;
  RECT 138.040 292.880 141.580 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER ME3 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER ME2 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER ME1 ;
  RECT 129.360 292.880 132.900 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER ME3 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER ME2 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER ME1 ;
  RECT 120.680 292.880 124.220 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER ME3 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER ME2 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER ME1 ;
  RECT 112.000 292.880 115.540 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER ME3 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER ME2 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER ME1 ;
  RECT 103.320 292.880 106.860 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER ME3 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER ME2 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER ME1 ;
  RECT 94.640 292.880 98.180 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER ME3 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER ME2 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER ME1 ;
  RECT 51.240 292.880 54.780 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER ME3 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER ME2 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER ME1 ;
  RECT 42.560 292.880 46.100 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER ME3 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER ME2 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER ME1 ;
  RECT 33.880 292.880 37.420 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER ME3 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER ME2 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER ME1 ;
  RECT 25.200 292.880 28.740 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER ME3 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER ME2 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER ME1 ;
  RECT 16.520 292.880 20.060 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER ME3 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER ME2 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER ME1 ;
  RECT 7.840 292.880 11.380 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER ME3 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER ME2 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER ME1 ;
  RECT 541.660 0.000 545.200 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER ME3 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER ME2 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER ME1 ;
  RECT 519.960 0.000 523.500 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER ME3 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER ME2 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER ME1 ;
  RECT 503.220 0.000 506.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER ME3 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER ME2 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER ME1 ;
  RECT 476.560 0.000 480.100 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.080 0.000 353.620 1.120 ;
  LAYER ME3 ;
  RECT 350.080 0.000 353.620 1.120 ;
  LAYER ME2 ;
  RECT 350.080 0.000 353.620 1.120 ;
  LAYER ME1 ;
  RECT 350.080 0.000 353.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.960 0.000 337.500 1.120 ;
  LAYER ME3 ;
  RECT 333.960 0.000 337.500 1.120 ;
  LAYER ME2 ;
  RECT 333.960 0.000 337.500 1.120 ;
  LAYER ME1 ;
  RECT 333.960 0.000 337.500 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER ME3 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER ME2 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER ME1 ;
  RECT 297.380 0.000 300.920 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 288.700 0.000 292.240 1.120 ;
  LAYER ME3 ;
  RECT 288.700 0.000 292.240 1.120 ;
  LAYER ME2 ;
  RECT 288.700 0.000 292.240 1.120 ;
  LAYER ME1 ;
  RECT 288.700 0.000 292.240 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER ME3 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER ME2 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER ME1 ;
  RECT 267.620 0.000 271.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME3 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME2 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME1 ;
  RECT 246.540 0.000 250.080 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER ME3 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER ME2 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER ME1 ;
  RECT 148.580 0.000 152.120 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 551.920 278.660 553.040 281.900 ;
  LAYER ME3 ;
  RECT 551.920 278.660 553.040 281.900 ;
  LAYER ME2 ;
  RECT 551.920 278.660 553.040 281.900 ;
  LAYER ME1 ;
  RECT 551.920 278.660 553.040 281.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 270.820 553.040 274.060 ;
  LAYER ME3 ;
  RECT 551.920 270.820 553.040 274.060 ;
  LAYER ME2 ;
  RECT 551.920 270.820 553.040 274.060 ;
  LAYER ME1 ;
  RECT 551.920 270.820 553.040 274.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 262.980 553.040 266.220 ;
  LAYER ME3 ;
  RECT 551.920 262.980 553.040 266.220 ;
  LAYER ME2 ;
  RECT 551.920 262.980 553.040 266.220 ;
  LAYER ME1 ;
  RECT 551.920 262.980 553.040 266.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 255.140 553.040 258.380 ;
  LAYER ME3 ;
  RECT 551.920 255.140 553.040 258.380 ;
  LAYER ME2 ;
  RECT 551.920 255.140 553.040 258.380 ;
  LAYER ME1 ;
  RECT 551.920 255.140 553.040 258.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 247.300 553.040 250.540 ;
  LAYER ME3 ;
  RECT 551.920 247.300 553.040 250.540 ;
  LAYER ME2 ;
  RECT 551.920 247.300 553.040 250.540 ;
  LAYER ME1 ;
  RECT 551.920 247.300 553.040 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 208.100 553.040 211.340 ;
  LAYER ME3 ;
  RECT 551.920 208.100 553.040 211.340 ;
  LAYER ME2 ;
  RECT 551.920 208.100 553.040 211.340 ;
  LAYER ME1 ;
  RECT 551.920 208.100 553.040 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 200.260 553.040 203.500 ;
  LAYER ME3 ;
  RECT 551.920 200.260 553.040 203.500 ;
  LAYER ME2 ;
  RECT 551.920 200.260 553.040 203.500 ;
  LAYER ME1 ;
  RECT 551.920 200.260 553.040 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 192.420 553.040 195.660 ;
  LAYER ME3 ;
  RECT 551.920 192.420 553.040 195.660 ;
  LAYER ME2 ;
  RECT 551.920 192.420 553.040 195.660 ;
  LAYER ME1 ;
  RECT 551.920 192.420 553.040 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 184.580 553.040 187.820 ;
  LAYER ME3 ;
  RECT 551.920 184.580 553.040 187.820 ;
  LAYER ME2 ;
  RECT 551.920 184.580 553.040 187.820 ;
  LAYER ME1 ;
  RECT 551.920 184.580 553.040 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 176.740 553.040 179.980 ;
  LAYER ME3 ;
  RECT 551.920 176.740 553.040 179.980 ;
  LAYER ME2 ;
  RECT 551.920 176.740 553.040 179.980 ;
  LAYER ME1 ;
  RECT 551.920 176.740 553.040 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 168.900 553.040 172.140 ;
  LAYER ME3 ;
  RECT 551.920 168.900 553.040 172.140 ;
  LAYER ME2 ;
  RECT 551.920 168.900 553.040 172.140 ;
  LAYER ME1 ;
  RECT 551.920 168.900 553.040 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 129.700 553.040 132.940 ;
  LAYER ME3 ;
  RECT 551.920 129.700 553.040 132.940 ;
  LAYER ME2 ;
  RECT 551.920 129.700 553.040 132.940 ;
  LAYER ME1 ;
  RECT 551.920 129.700 553.040 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 121.860 553.040 125.100 ;
  LAYER ME3 ;
  RECT 551.920 121.860 553.040 125.100 ;
  LAYER ME2 ;
  RECT 551.920 121.860 553.040 125.100 ;
  LAYER ME1 ;
  RECT 551.920 121.860 553.040 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 114.020 553.040 117.260 ;
  LAYER ME3 ;
  RECT 551.920 114.020 553.040 117.260 ;
  LAYER ME2 ;
  RECT 551.920 114.020 553.040 117.260 ;
  LAYER ME1 ;
  RECT 551.920 114.020 553.040 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 106.180 553.040 109.420 ;
  LAYER ME3 ;
  RECT 551.920 106.180 553.040 109.420 ;
  LAYER ME2 ;
  RECT 551.920 106.180 553.040 109.420 ;
  LAYER ME1 ;
  RECT 551.920 106.180 553.040 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 98.340 553.040 101.580 ;
  LAYER ME3 ;
  RECT 551.920 98.340 553.040 101.580 ;
  LAYER ME2 ;
  RECT 551.920 98.340 553.040 101.580 ;
  LAYER ME1 ;
  RECT 551.920 98.340 553.040 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 90.500 553.040 93.740 ;
  LAYER ME3 ;
  RECT 551.920 90.500 553.040 93.740 ;
  LAYER ME2 ;
  RECT 551.920 90.500 553.040 93.740 ;
  LAYER ME1 ;
  RECT 551.920 90.500 553.040 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 51.300 553.040 54.540 ;
  LAYER ME3 ;
  RECT 551.920 51.300 553.040 54.540 ;
  LAYER ME2 ;
  RECT 551.920 51.300 553.040 54.540 ;
  LAYER ME1 ;
  RECT 551.920 51.300 553.040 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 43.460 553.040 46.700 ;
  LAYER ME3 ;
  RECT 551.920 43.460 553.040 46.700 ;
  LAYER ME2 ;
  RECT 551.920 43.460 553.040 46.700 ;
  LAYER ME1 ;
  RECT 551.920 43.460 553.040 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 35.620 553.040 38.860 ;
  LAYER ME3 ;
  RECT 551.920 35.620 553.040 38.860 ;
  LAYER ME2 ;
  RECT 551.920 35.620 553.040 38.860 ;
  LAYER ME1 ;
  RECT 551.920 35.620 553.040 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 27.780 553.040 31.020 ;
  LAYER ME3 ;
  RECT 551.920 27.780 553.040 31.020 ;
  LAYER ME2 ;
  RECT 551.920 27.780 553.040 31.020 ;
  LAYER ME1 ;
  RECT 551.920 27.780 553.040 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 19.940 553.040 23.180 ;
  LAYER ME3 ;
  RECT 551.920 19.940 553.040 23.180 ;
  LAYER ME2 ;
  RECT 551.920 19.940 553.040 23.180 ;
  LAYER ME1 ;
  RECT 551.920 19.940 553.040 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.920 12.100 553.040 15.340 ;
  LAYER ME3 ;
  RECT 551.920 12.100 553.040 15.340 ;
  LAYER ME2 ;
  RECT 551.920 12.100 553.040 15.340 ;
  LAYER ME1 ;
  RECT 551.920 12.100 553.040 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.660 292.880 545.200 294.000 ;
  LAYER ME3 ;
  RECT 541.660 292.880 545.200 294.000 ;
  LAYER ME2 ;
  RECT 541.660 292.880 545.200 294.000 ;
  LAYER ME1 ;
  RECT 541.660 292.880 545.200 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.980 292.880 536.520 294.000 ;
  LAYER ME3 ;
  RECT 532.980 292.880 536.520 294.000 ;
  LAYER ME2 ;
  RECT 532.980 292.880 536.520 294.000 ;
  LAYER ME1 ;
  RECT 532.980 292.880 536.520 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.580 292.880 493.120 294.000 ;
  LAYER ME3 ;
  RECT 489.580 292.880 493.120 294.000 ;
  LAYER ME2 ;
  RECT 489.580 292.880 493.120 294.000 ;
  LAYER ME1 ;
  RECT 489.580 292.880 493.120 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.900 292.880 484.440 294.000 ;
  LAYER ME3 ;
  RECT 480.900 292.880 484.440 294.000 ;
  LAYER ME2 ;
  RECT 480.900 292.880 484.440 294.000 ;
  LAYER ME1 ;
  RECT 480.900 292.880 484.440 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 292.880 475.760 294.000 ;
  LAYER ME3 ;
  RECT 472.220 292.880 475.760 294.000 ;
  LAYER ME2 ;
  RECT 472.220 292.880 475.760 294.000 ;
  LAYER ME1 ;
  RECT 472.220 292.880 475.760 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.540 292.880 467.080 294.000 ;
  LAYER ME3 ;
  RECT 463.540 292.880 467.080 294.000 ;
  LAYER ME2 ;
  RECT 463.540 292.880 467.080 294.000 ;
  LAYER ME1 ;
  RECT 463.540 292.880 467.080 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.860 292.880 458.400 294.000 ;
  LAYER ME3 ;
  RECT 454.860 292.880 458.400 294.000 ;
  LAYER ME2 ;
  RECT 454.860 292.880 458.400 294.000 ;
  LAYER ME1 ;
  RECT 454.860 292.880 458.400 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.180 292.880 449.720 294.000 ;
  LAYER ME3 ;
  RECT 446.180 292.880 449.720 294.000 ;
  LAYER ME2 ;
  RECT 446.180 292.880 449.720 294.000 ;
  LAYER ME1 ;
  RECT 446.180 292.880 449.720 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 292.880 406.320 294.000 ;
  LAYER ME3 ;
  RECT 402.780 292.880 406.320 294.000 ;
  LAYER ME2 ;
  RECT 402.780 292.880 406.320 294.000 ;
  LAYER ME1 ;
  RECT 402.780 292.880 406.320 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.100 292.880 397.640 294.000 ;
  LAYER ME3 ;
  RECT 394.100 292.880 397.640 294.000 ;
  LAYER ME2 ;
  RECT 394.100 292.880 397.640 294.000 ;
  LAYER ME1 ;
  RECT 394.100 292.880 397.640 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.420 292.880 388.960 294.000 ;
  LAYER ME3 ;
  RECT 385.420 292.880 388.960 294.000 ;
  LAYER ME2 ;
  RECT 385.420 292.880 388.960 294.000 ;
  LAYER ME1 ;
  RECT 385.420 292.880 388.960 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.740 292.880 380.280 294.000 ;
  LAYER ME3 ;
  RECT 376.740 292.880 380.280 294.000 ;
  LAYER ME2 ;
  RECT 376.740 292.880 380.280 294.000 ;
  LAYER ME1 ;
  RECT 376.740 292.880 380.280 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.060 292.880 371.600 294.000 ;
  LAYER ME3 ;
  RECT 368.060 292.880 371.600 294.000 ;
  LAYER ME2 ;
  RECT 368.060 292.880 371.600 294.000 ;
  LAYER ME1 ;
  RECT 368.060 292.880 371.600 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.380 292.880 362.920 294.000 ;
  LAYER ME3 ;
  RECT 359.380 292.880 362.920 294.000 ;
  LAYER ME2 ;
  RECT 359.380 292.880 362.920 294.000 ;
  LAYER ME1 ;
  RECT 359.380 292.880 362.920 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.980 292.880 319.520 294.000 ;
  LAYER ME3 ;
  RECT 315.980 292.880 319.520 294.000 ;
  LAYER ME2 ;
  RECT 315.980 292.880 319.520 294.000 ;
  LAYER ME1 ;
  RECT 315.980 292.880 319.520 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER ME3 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER ME2 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER ME1 ;
  RECT 307.300 292.880 310.840 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER ME3 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER ME2 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER ME1 ;
  RECT 298.620 292.880 302.160 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER ME3 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER ME2 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER ME1 ;
  RECT 289.940 292.880 293.480 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER ME3 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER ME2 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER ME1 ;
  RECT 281.260 292.880 284.800 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER ME3 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER ME2 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER ME1 ;
  RECT 272.580 292.880 276.120 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER ME3 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER ME2 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER ME1 ;
  RECT 229.180 292.880 232.720 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER ME3 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER ME2 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER ME1 ;
  RECT 220.500 292.880 224.040 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER ME3 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER ME2 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER ME1 ;
  RECT 211.820 292.880 215.360 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER ME3 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER ME2 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER ME1 ;
  RECT 203.140 292.880 206.680 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER ME3 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER ME2 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER ME1 ;
  RECT 194.460 292.880 198.000 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER ME3 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER ME2 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER ME1 ;
  RECT 185.780 292.880 189.320 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER ME3 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER ME2 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER ME1 ;
  RECT 142.380 292.880 145.920 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER ME3 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER ME2 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER ME1 ;
  RECT 133.700 292.880 137.240 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER ME3 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER ME2 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER ME1 ;
  RECT 125.020 292.880 128.560 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER ME3 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER ME2 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER ME1 ;
  RECT 116.340 292.880 119.880 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER ME3 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER ME2 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER ME1 ;
  RECT 107.660 292.880 111.200 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER ME3 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER ME2 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER ME1 ;
  RECT 98.980 292.880 102.520 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER ME3 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER ME2 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER ME1 ;
  RECT 55.580 292.880 59.120 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER ME3 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER ME2 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER ME1 ;
  RECT 46.900 292.880 50.440 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER ME3 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER ME2 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER ME1 ;
  RECT 38.220 292.880 41.760 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER ME3 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER ME2 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER ME1 ;
  RECT 29.540 292.880 33.080 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER ME3 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER ME2 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER ME1 ;
  RECT 20.860 292.880 24.400 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER ME3 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER ME2 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER ME1 ;
  RECT 12.180 292.880 15.720 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER ME3 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER ME2 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER ME1 ;
  RECT 532.980 0.000 536.520 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER ME3 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER ME2 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER ME1 ;
  RECT 511.900 0.000 515.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER ME3 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER ME2 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER ME1 ;
  RECT 490.200 0.000 493.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 0.000 367.260 1.120 ;
  LAYER ME3 ;
  RECT 363.720 0.000 367.260 1.120 ;
  LAYER ME2 ;
  RECT 363.720 0.000 367.260 1.120 ;
  LAYER ME1 ;
  RECT 363.720 0.000 367.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER ME3 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER ME2 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER ME1 ;
  RECT 342.020 0.000 345.560 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.920 0.000 311.460 1.120 ;
  LAYER ME3 ;
  RECT 307.920 0.000 311.460 1.120 ;
  LAYER ME2 ;
  RECT 307.920 0.000 311.460 1.120 ;
  LAYER ME1 ;
  RECT 307.920 0.000 311.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.040 0.000 296.580 1.120 ;
  LAYER ME3 ;
  RECT 293.040 0.000 296.580 1.120 ;
  LAYER ME2 ;
  RECT 293.040 0.000 296.580 1.120 ;
  LAYER ME1 ;
  RECT 293.040 0.000 296.580 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 284.360 0.000 287.900 1.120 ;
  LAYER ME3 ;
  RECT 284.360 0.000 287.900 1.120 ;
  LAYER ME2 ;
  RECT 284.360 0.000 287.900 1.120 ;
  LAYER ME1 ;
  RECT 284.360 0.000 287.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER ME3 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER ME2 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER ME1 ;
  RECT 257.080 0.000 260.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.640 0.000 160.180 1.120 ;
  LAYER ME3 ;
  RECT 156.640 0.000 160.180 1.120 ;
  LAYER ME2 ;
  RECT 156.640 0.000 160.180 1.120 ;
  LAYER ME1 ;
  RECT 156.640 0.000 160.180 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
END GND
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER ME3 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER ME2 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER ME1 ;
  RECT 539.460 0.000 540.580 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER ME3 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER ME2 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER ME1 ;
  RECT 530.780 0.000 531.900 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER ME3 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER ME2 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER ME1 ;
  RECT 525.820 0.000 526.940 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER ME3 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER ME2 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER ME1 ;
  RECT 517.760 0.000 518.880 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME3 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME2 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME1 ;
  RECT 509.700 0.000 510.820 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER ME3 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER ME2 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER ME1 ;
  RECT 501.020 0.000 502.140 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER ME3 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER ME2 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER ME1 ;
  RECT 496.060 0.000 497.180 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER ME3 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER ME2 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER ME1 ;
  RECT 483.040 0.000 484.160 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER ME3 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER ME2 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER ME1 ;
  RECT 474.360 0.000 475.480 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER ME3 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER ME2 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER ME1 ;
  RECT 469.400 0.000 470.520 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER ME3 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER ME2 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER ME1 ;
  RECT 461.340 0.000 462.460 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER ME3 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER ME2 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER ME1 ;
  RECT 452.660 0.000 453.780 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER ME3 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER ME2 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER ME1 ;
  RECT 444.600 0.000 445.720 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER ME3 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER ME2 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER ME1 ;
  RECT 439.640 0.000 440.760 1.120 ;
 END
END DO24
PIN WEB3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 435.300 0.000 436.420 1.120 ;
  LAYER ME3 ;
  RECT 435.300 0.000 436.420 1.120 ;
  LAYER ME2 ;
  RECT 435.300 0.000 436.420 1.120 ;
  LAYER ME1 ;
  RECT 435.300 0.000 436.420 1.120 ;
 END
END WEB3
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER ME3 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER ME2 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER ME1 ;
  RECT 430.960 0.000 432.080 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER ME3 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER ME2 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER ME1 ;
  RECT 426.620 0.000 427.740 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER ME3 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER ME2 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER ME1 ;
  RECT 417.940 0.000 419.060 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER ME3 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER ME2 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER ME1 ;
  RECT 412.980 0.000 414.100 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER ME3 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER ME2 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER ME1 ;
  RECT 404.920 0.000 406.040 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER ME3 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER ME2 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER ME1 ;
  RECT 396.240 0.000 397.360 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 388.180 0.000 389.300 1.120 ;
  LAYER ME3 ;
  RECT 388.180 0.000 389.300 1.120 ;
  LAYER ME2 ;
  RECT 388.180 0.000 389.300 1.120 ;
  LAYER ME1 ;
  RECT 388.180 0.000 389.300 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER ME3 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER ME2 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER ME1 ;
  RECT 383.220 0.000 384.340 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER ME3 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER ME2 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER ME1 ;
  RECT 374.540 0.000 375.660 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 369.580 0.000 370.700 1.120 ;
  LAYER ME3 ;
  RECT 369.580 0.000 370.700 1.120 ;
  LAYER ME2 ;
  RECT 369.580 0.000 370.700 1.120 ;
  LAYER ME1 ;
  RECT 369.580 0.000 370.700 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 361.520 0.000 362.640 1.120 ;
  LAYER ME3 ;
  RECT 361.520 0.000 362.640 1.120 ;
  LAYER ME2 ;
  RECT 361.520 0.000 362.640 1.120 ;
  LAYER ME1 ;
  RECT 361.520 0.000 362.640 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER ME3 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER ME2 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER ME1 ;
  RECT 356.560 0.000 357.680 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 347.880 0.000 349.000 1.120 ;
  LAYER ME3 ;
  RECT 347.880 0.000 349.000 1.120 ;
  LAYER ME2 ;
  RECT 347.880 0.000 349.000 1.120 ;
  LAYER ME1 ;
  RECT 347.880 0.000 349.000 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 339.820 0.000 340.940 1.120 ;
  LAYER ME3 ;
  RECT 339.820 0.000 340.940 1.120 ;
  LAYER ME2 ;
  RECT 339.820 0.000 340.940 1.120 ;
  LAYER ME1 ;
  RECT 339.820 0.000 340.940 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 331.760 0.000 332.880 1.120 ;
  LAYER ME3 ;
  RECT 331.760 0.000 332.880 1.120 ;
  LAYER ME2 ;
  RECT 331.760 0.000 332.880 1.120 ;
  LAYER ME1 ;
  RECT 331.760 0.000 332.880 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER ME3 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER ME2 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER ME1 ;
  RECT 326.800 0.000 327.920 1.120 ;
 END
END DO16
PIN WEB2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER ME3 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER ME2 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER ME1 ;
  RECT 321.840 0.000 322.960 1.120 ;
 END
END WEB2
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 318.120 0.000 319.240 1.120 ;
  LAYER ME3 ;
  RECT 318.120 0.000 319.240 1.120 ;
  LAYER ME2 ;
  RECT 318.120 0.000 319.240 1.120 ;
  LAYER ME1 ;
  RECT 318.120 0.000 319.240 1.120 ;
 END
END DI16
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 312.540 0.000 313.660 1.120 ;
  LAYER ME3 ;
  RECT 312.540 0.000 313.660 1.120 ;
  LAYER ME2 ;
  RECT 312.540 0.000 313.660 1.120 ;
  LAYER ME1 ;
  RECT 312.540 0.000 313.660 1.120 ;
 END
END A1
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 305.720 0.000 306.840 1.120 ;
  LAYER ME3 ;
  RECT 305.720 0.000 306.840 1.120 ;
  LAYER ME2 ;
  RECT 305.720 0.000 306.840 1.120 ;
  LAYER ME1 ;
  RECT 305.720 0.000 306.840 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 303.860 0.000 304.980 1.120 ;
  LAYER ME3 ;
  RECT 303.860 0.000 304.980 1.120 ;
  LAYER ME2 ;
  RECT 303.860 0.000 304.980 1.120 ;
  LAYER ME1 ;
  RECT 303.860 0.000 304.980 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER ME3 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER ME2 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER ME1 ;
  RECT 282.160 0.000 283.280 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER ME3 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER ME2 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER ME1 ;
  RECT 279.060 0.000 280.180 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 277.200 0.000 278.320 1.120 ;
  LAYER ME3 ;
  RECT 277.200 0.000 278.320 1.120 ;
  LAYER ME2 ;
  RECT 277.200 0.000 278.320 1.120 ;
  LAYER ME1 ;
  RECT 277.200 0.000 278.320 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER ME3 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER ME2 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER ME1 ;
  RECT 272.860 0.000 273.980 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER ME3 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER ME2 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER ME1 ;
  RECT 265.420 0.000 266.540 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME3 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME2 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME1 ;
  RECT 262.320 0.000 263.440 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME3 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME2 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME1 ;
  RECT 251.780 0.000 252.900 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME3 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME2 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME1 ;
  RECT 244.340 0.000 245.460 1.120 ;
 END
END A8
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN WEB1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 128.400 0.000 129.520 1.120 ;
  LAYER ME3 ;
  RECT 128.400 0.000 129.520 1.120 ;
  LAYER ME2 ;
  RECT 128.400 0.000 129.520 1.120 ;
  LAYER ME1 ;
  RECT 128.400 0.000 129.520 1.120 ;
 END
END WEB1
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN WEB0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER ME3 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER ME2 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER ME1 ;
  RECT 15.560 0.000 16.680 1.120 ;
 END
END WEB0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 553.040 294.000 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 553.040 294.000 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 553.040 294.000 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 553.040 294.000 ;
  LAYER VI1 ;
  RECT 0.000 0.140 553.040 294.000 ;
  LAYER VI2 ;
  RECT 0.000 0.140 553.040 294.000 ;
  LAYER VI3 ;
  RECT 0.000 0.140 553.040 294.000 ;
END
END SRAM_small
END LIBRARY



