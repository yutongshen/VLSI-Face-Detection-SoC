PLIC/PLIC.sv