../include/AHB_def.svh