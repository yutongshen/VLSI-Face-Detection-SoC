AHB/AHB.sv