../include/ALUCtrl.svh