AHB/MuxS2M.sv