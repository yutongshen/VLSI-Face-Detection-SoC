parameter [2:0] FUNCT3_ADD_SUB   = 3'b000,
                FUNCT3_SLL       = 3'b001,
                FUNCT3_SLT       = 3'b010,
                FUNCT3_SLTU      = 3'b011,
                FUNCT3_XOR       = 3'b100,
                FUNCT3_SRL_SRA   = 3'b101,
                FUNCT3_OR        = 3'b110,
                FUNCT3_AND       = 3'b111,

                FUNCT3_ADDI_JALR = 3'b000,
                FUNCT3_SLLI      = 3'b001,
                FUNCT3_SLTI      = 3'b010,
                FUNCT3_SLTIU     = 3'b011,
                FUNCT3_XORI      = 3'b100,
                FUNCT3_SRLI_SRAI = 3'b101,
                FUNCT3_ORI       = 3'b110,
                FUNCT3_ANDI      = 3'b111,

                FUNCT3_BEQ       = 3'b000,
                FUNCT3_BNE       = 3'b001,
                FUNCT3_BLT       = 3'b100,
                FUNCT3_BGE       = 3'b101,
                FUNCT3_BLTU      = 3'b110,
                FUNCT3_BGEU      = 3'b111;
