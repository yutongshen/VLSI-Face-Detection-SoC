# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SUMA180_8192X8X4BM2
#       Words            : 8192
#       Bits             : 8
#       Byte-Write       : 4
#       Aspect Ratio     : 2
#       Output Loading   : 0.01  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2019/01/15 02:45:38
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SUMA180_8192X8X4BM2
CLASS BLOCK ;
FOREIGN SUMA180_8192X8X4BM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 1015.560 BY 1391.600 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 1014.440 1380.180 1015.560 1383.420 ;
  LAYER ME3 ;
  RECT 1014.440 1380.180 1015.560 1383.420 ;
  LAYER ME2 ;
  RECT 1014.440 1380.180 1015.560 1383.420 ;
  LAYER ME1 ;
  RECT 1014.440 1380.180 1015.560 1383.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1372.340 1015.560 1375.580 ;
  LAYER ME3 ;
  RECT 1014.440 1372.340 1015.560 1375.580 ;
  LAYER ME2 ;
  RECT 1014.440 1372.340 1015.560 1375.580 ;
  LAYER ME1 ;
  RECT 1014.440 1372.340 1015.560 1375.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1364.500 1015.560 1367.740 ;
  LAYER ME3 ;
  RECT 1014.440 1364.500 1015.560 1367.740 ;
  LAYER ME2 ;
  RECT 1014.440 1364.500 1015.560 1367.740 ;
  LAYER ME1 ;
  RECT 1014.440 1364.500 1015.560 1367.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1356.660 1015.560 1359.900 ;
  LAYER ME3 ;
  RECT 1014.440 1356.660 1015.560 1359.900 ;
  LAYER ME2 ;
  RECT 1014.440 1356.660 1015.560 1359.900 ;
  LAYER ME1 ;
  RECT 1014.440 1356.660 1015.560 1359.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1348.820 1015.560 1352.060 ;
  LAYER ME3 ;
  RECT 1014.440 1348.820 1015.560 1352.060 ;
  LAYER ME2 ;
  RECT 1014.440 1348.820 1015.560 1352.060 ;
  LAYER ME1 ;
  RECT 1014.440 1348.820 1015.560 1352.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1340.980 1015.560 1344.220 ;
  LAYER ME3 ;
  RECT 1014.440 1340.980 1015.560 1344.220 ;
  LAYER ME2 ;
  RECT 1014.440 1340.980 1015.560 1344.220 ;
  LAYER ME1 ;
  RECT 1014.440 1340.980 1015.560 1344.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1301.780 1015.560 1305.020 ;
  LAYER ME3 ;
  RECT 1014.440 1301.780 1015.560 1305.020 ;
  LAYER ME2 ;
  RECT 1014.440 1301.780 1015.560 1305.020 ;
  LAYER ME1 ;
  RECT 1014.440 1301.780 1015.560 1305.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1293.940 1015.560 1297.180 ;
  LAYER ME3 ;
  RECT 1014.440 1293.940 1015.560 1297.180 ;
  LAYER ME2 ;
  RECT 1014.440 1293.940 1015.560 1297.180 ;
  LAYER ME1 ;
  RECT 1014.440 1293.940 1015.560 1297.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1286.100 1015.560 1289.340 ;
  LAYER ME3 ;
  RECT 1014.440 1286.100 1015.560 1289.340 ;
  LAYER ME2 ;
  RECT 1014.440 1286.100 1015.560 1289.340 ;
  LAYER ME1 ;
  RECT 1014.440 1286.100 1015.560 1289.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1278.260 1015.560 1281.500 ;
  LAYER ME3 ;
  RECT 1014.440 1278.260 1015.560 1281.500 ;
  LAYER ME2 ;
  RECT 1014.440 1278.260 1015.560 1281.500 ;
  LAYER ME1 ;
  RECT 1014.440 1278.260 1015.560 1281.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1270.420 1015.560 1273.660 ;
  LAYER ME3 ;
  RECT 1014.440 1270.420 1015.560 1273.660 ;
  LAYER ME2 ;
  RECT 1014.440 1270.420 1015.560 1273.660 ;
  LAYER ME1 ;
  RECT 1014.440 1270.420 1015.560 1273.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1262.580 1015.560 1265.820 ;
  LAYER ME3 ;
  RECT 1014.440 1262.580 1015.560 1265.820 ;
  LAYER ME2 ;
  RECT 1014.440 1262.580 1015.560 1265.820 ;
  LAYER ME1 ;
  RECT 1014.440 1262.580 1015.560 1265.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1223.380 1015.560 1226.620 ;
  LAYER ME3 ;
  RECT 1014.440 1223.380 1015.560 1226.620 ;
  LAYER ME2 ;
  RECT 1014.440 1223.380 1015.560 1226.620 ;
  LAYER ME1 ;
  RECT 1014.440 1223.380 1015.560 1226.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1215.540 1015.560 1218.780 ;
  LAYER ME3 ;
  RECT 1014.440 1215.540 1015.560 1218.780 ;
  LAYER ME2 ;
  RECT 1014.440 1215.540 1015.560 1218.780 ;
  LAYER ME1 ;
  RECT 1014.440 1215.540 1015.560 1218.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1207.700 1015.560 1210.940 ;
  LAYER ME3 ;
  RECT 1014.440 1207.700 1015.560 1210.940 ;
  LAYER ME2 ;
  RECT 1014.440 1207.700 1015.560 1210.940 ;
  LAYER ME1 ;
  RECT 1014.440 1207.700 1015.560 1210.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1199.860 1015.560 1203.100 ;
  LAYER ME3 ;
  RECT 1014.440 1199.860 1015.560 1203.100 ;
  LAYER ME2 ;
  RECT 1014.440 1199.860 1015.560 1203.100 ;
  LAYER ME1 ;
  RECT 1014.440 1199.860 1015.560 1203.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1192.020 1015.560 1195.260 ;
  LAYER ME3 ;
  RECT 1014.440 1192.020 1015.560 1195.260 ;
  LAYER ME2 ;
  RECT 1014.440 1192.020 1015.560 1195.260 ;
  LAYER ME1 ;
  RECT 1014.440 1192.020 1015.560 1195.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1184.180 1015.560 1187.420 ;
  LAYER ME3 ;
  RECT 1014.440 1184.180 1015.560 1187.420 ;
  LAYER ME2 ;
  RECT 1014.440 1184.180 1015.560 1187.420 ;
  LAYER ME1 ;
  RECT 1014.440 1184.180 1015.560 1187.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1144.980 1015.560 1148.220 ;
  LAYER ME3 ;
  RECT 1014.440 1144.980 1015.560 1148.220 ;
  LAYER ME2 ;
  RECT 1014.440 1144.980 1015.560 1148.220 ;
  LAYER ME1 ;
  RECT 1014.440 1144.980 1015.560 1148.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1137.140 1015.560 1140.380 ;
  LAYER ME3 ;
  RECT 1014.440 1137.140 1015.560 1140.380 ;
  LAYER ME2 ;
  RECT 1014.440 1137.140 1015.560 1140.380 ;
  LAYER ME1 ;
  RECT 1014.440 1137.140 1015.560 1140.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1129.300 1015.560 1132.540 ;
  LAYER ME3 ;
  RECT 1014.440 1129.300 1015.560 1132.540 ;
  LAYER ME2 ;
  RECT 1014.440 1129.300 1015.560 1132.540 ;
  LAYER ME1 ;
  RECT 1014.440 1129.300 1015.560 1132.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1121.460 1015.560 1124.700 ;
  LAYER ME3 ;
  RECT 1014.440 1121.460 1015.560 1124.700 ;
  LAYER ME2 ;
  RECT 1014.440 1121.460 1015.560 1124.700 ;
  LAYER ME1 ;
  RECT 1014.440 1121.460 1015.560 1124.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1113.620 1015.560 1116.860 ;
  LAYER ME3 ;
  RECT 1014.440 1113.620 1015.560 1116.860 ;
  LAYER ME2 ;
  RECT 1014.440 1113.620 1015.560 1116.860 ;
  LAYER ME1 ;
  RECT 1014.440 1113.620 1015.560 1116.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1105.780 1015.560 1109.020 ;
  LAYER ME3 ;
  RECT 1014.440 1105.780 1015.560 1109.020 ;
  LAYER ME2 ;
  RECT 1014.440 1105.780 1015.560 1109.020 ;
  LAYER ME1 ;
  RECT 1014.440 1105.780 1015.560 1109.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1066.580 1015.560 1069.820 ;
  LAYER ME3 ;
  RECT 1014.440 1066.580 1015.560 1069.820 ;
  LAYER ME2 ;
  RECT 1014.440 1066.580 1015.560 1069.820 ;
  LAYER ME1 ;
  RECT 1014.440 1066.580 1015.560 1069.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1058.740 1015.560 1061.980 ;
  LAYER ME3 ;
  RECT 1014.440 1058.740 1015.560 1061.980 ;
  LAYER ME2 ;
  RECT 1014.440 1058.740 1015.560 1061.980 ;
  LAYER ME1 ;
  RECT 1014.440 1058.740 1015.560 1061.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1050.900 1015.560 1054.140 ;
  LAYER ME3 ;
  RECT 1014.440 1050.900 1015.560 1054.140 ;
  LAYER ME2 ;
  RECT 1014.440 1050.900 1015.560 1054.140 ;
  LAYER ME1 ;
  RECT 1014.440 1050.900 1015.560 1054.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1043.060 1015.560 1046.300 ;
  LAYER ME3 ;
  RECT 1014.440 1043.060 1015.560 1046.300 ;
  LAYER ME2 ;
  RECT 1014.440 1043.060 1015.560 1046.300 ;
  LAYER ME1 ;
  RECT 1014.440 1043.060 1015.560 1046.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1035.220 1015.560 1038.460 ;
  LAYER ME3 ;
  RECT 1014.440 1035.220 1015.560 1038.460 ;
  LAYER ME2 ;
  RECT 1014.440 1035.220 1015.560 1038.460 ;
  LAYER ME1 ;
  RECT 1014.440 1035.220 1015.560 1038.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1027.380 1015.560 1030.620 ;
  LAYER ME3 ;
  RECT 1014.440 1027.380 1015.560 1030.620 ;
  LAYER ME2 ;
  RECT 1014.440 1027.380 1015.560 1030.620 ;
  LAYER ME1 ;
  RECT 1014.440 1027.380 1015.560 1030.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 988.180 1015.560 991.420 ;
  LAYER ME3 ;
  RECT 1014.440 988.180 1015.560 991.420 ;
  LAYER ME2 ;
  RECT 1014.440 988.180 1015.560 991.420 ;
  LAYER ME1 ;
  RECT 1014.440 988.180 1015.560 991.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 980.340 1015.560 983.580 ;
  LAYER ME3 ;
  RECT 1014.440 980.340 1015.560 983.580 ;
  LAYER ME2 ;
  RECT 1014.440 980.340 1015.560 983.580 ;
  LAYER ME1 ;
  RECT 1014.440 980.340 1015.560 983.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 972.500 1015.560 975.740 ;
  LAYER ME3 ;
  RECT 1014.440 972.500 1015.560 975.740 ;
  LAYER ME2 ;
  RECT 1014.440 972.500 1015.560 975.740 ;
  LAYER ME1 ;
  RECT 1014.440 972.500 1015.560 975.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 964.660 1015.560 967.900 ;
  LAYER ME3 ;
  RECT 1014.440 964.660 1015.560 967.900 ;
  LAYER ME2 ;
  RECT 1014.440 964.660 1015.560 967.900 ;
  LAYER ME1 ;
  RECT 1014.440 964.660 1015.560 967.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 956.820 1015.560 960.060 ;
  LAYER ME3 ;
  RECT 1014.440 956.820 1015.560 960.060 ;
  LAYER ME2 ;
  RECT 1014.440 956.820 1015.560 960.060 ;
  LAYER ME1 ;
  RECT 1014.440 956.820 1015.560 960.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 948.980 1015.560 952.220 ;
  LAYER ME3 ;
  RECT 1014.440 948.980 1015.560 952.220 ;
  LAYER ME2 ;
  RECT 1014.440 948.980 1015.560 952.220 ;
  LAYER ME1 ;
  RECT 1014.440 948.980 1015.560 952.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 909.780 1015.560 913.020 ;
  LAYER ME3 ;
  RECT 1014.440 909.780 1015.560 913.020 ;
  LAYER ME2 ;
  RECT 1014.440 909.780 1015.560 913.020 ;
  LAYER ME1 ;
  RECT 1014.440 909.780 1015.560 913.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 901.940 1015.560 905.180 ;
  LAYER ME3 ;
  RECT 1014.440 901.940 1015.560 905.180 ;
  LAYER ME2 ;
  RECT 1014.440 901.940 1015.560 905.180 ;
  LAYER ME1 ;
  RECT 1014.440 901.940 1015.560 905.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 894.100 1015.560 897.340 ;
  LAYER ME3 ;
  RECT 1014.440 894.100 1015.560 897.340 ;
  LAYER ME2 ;
  RECT 1014.440 894.100 1015.560 897.340 ;
  LAYER ME1 ;
  RECT 1014.440 894.100 1015.560 897.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 886.260 1015.560 889.500 ;
  LAYER ME3 ;
  RECT 1014.440 886.260 1015.560 889.500 ;
  LAYER ME2 ;
  RECT 1014.440 886.260 1015.560 889.500 ;
  LAYER ME1 ;
  RECT 1014.440 886.260 1015.560 889.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 878.420 1015.560 881.660 ;
  LAYER ME3 ;
  RECT 1014.440 878.420 1015.560 881.660 ;
  LAYER ME2 ;
  RECT 1014.440 878.420 1015.560 881.660 ;
  LAYER ME1 ;
  RECT 1014.440 878.420 1015.560 881.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 870.580 1015.560 873.820 ;
  LAYER ME3 ;
  RECT 1014.440 870.580 1015.560 873.820 ;
  LAYER ME2 ;
  RECT 1014.440 870.580 1015.560 873.820 ;
  LAYER ME1 ;
  RECT 1014.440 870.580 1015.560 873.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 831.380 1015.560 834.620 ;
  LAYER ME3 ;
  RECT 1014.440 831.380 1015.560 834.620 ;
  LAYER ME2 ;
  RECT 1014.440 831.380 1015.560 834.620 ;
  LAYER ME1 ;
  RECT 1014.440 831.380 1015.560 834.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 823.540 1015.560 826.780 ;
  LAYER ME3 ;
  RECT 1014.440 823.540 1015.560 826.780 ;
  LAYER ME2 ;
  RECT 1014.440 823.540 1015.560 826.780 ;
  LAYER ME1 ;
  RECT 1014.440 823.540 1015.560 826.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 815.700 1015.560 818.940 ;
  LAYER ME3 ;
  RECT 1014.440 815.700 1015.560 818.940 ;
  LAYER ME2 ;
  RECT 1014.440 815.700 1015.560 818.940 ;
  LAYER ME1 ;
  RECT 1014.440 815.700 1015.560 818.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 807.860 1015.560 811.100 ;
  LAYER ME3 ;
  RECT 1014.440 807.860 1015.560 811.100 ;
  LAYER ME2 ;
  RECT 1014.440 807.860 1015.560 811.100 ;
  LAYER ME1 ;
  RECT 1014.440 807.860 1015.560 811.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 800.020 1015.560 803.260 ;
  LAYER ME3 ;
  RECT 1014.440 800.020 1015.560 803.260 ;
  LAYER ME2 ;
  RECT 1014.440 800.020 1015.560 803.260 ;
  LAYER ME1 ;
  RECT 1014.440 800.020 1015.560 803.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 792.180 1015.560 795.420 ;
  LAYER ME3 ;
  RECT 1014.440 792.180 1015.560 795.420 ;
  LAYER ME2 ;
  RECT 1014.440 792.180 1015.560 795.420 ;
  LAYER ME1 ;
  RECT 1014.440 792.180 1015.560 795.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 752.980 1015.560 756.220 ;
  LAYER ME3 ;
  RECT 1014.440 752.980 1015.560 756.220 ;
  LAYER ME2 ;
  RECT 1014.440 752.980 1015.560 756.220 ;
  LAYER ME1 ;
  RECT 1014.440 752.980 1015.560 756.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 745.140 1015.560 748.380 ;
  LAYER ME3 ;
  RECT 1014.440 745.140 1015.560 748.380 ;
  LAYER ME2 ;
  RECT 1014.440 745.140 1015.560 748.380 ;
  LAYER ME1 ;
  RECT 1014.440 745.140 1015.560 748.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 737.300 1015.560 740.540 ;
  LAYER ME3 ;
  RECT 1014.440 737.300 1015.560 740.540 ;
  LAYER ME2 ;
  RECT 1014.440 737.300 1015.560 740.540 ;
  LAYER ME1 ;
  RECT 1014.440 737.300 1015.560 740.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 729.460 1015.560 732.700 ;
  LAYER ME3 ;
  RECT 1014.440 729.460 1015.560 732.700 ;
  LAYER ME2 ;
  RECT 1014.440 729.460 1015.560 732.700 ;
  LAYER ME1 ;
  RECT 1014.440 729.460 1015.560 732.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 721.620 1015.560 724.860 ;
  LAYER ME3 ;
  RECT 1014.440 721.620 1015.560 724.860 ;
  LAYER ME2 ;
  RECT 1014.440 721.620 1015.560 724.860 ;
  LAYER ME1 ;
  RECT 1014.440 721.620 1015.560 724.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 713.780 1015.560 717.020 ;
  LAYER ME3 ;
  RECT 1014.440 713.780 1015.560 717.020 ;
  LAYER ME2 ;
  RECT 1014.440 713.780 1015.560 717.020 ;
  LAYER ME1 ;
  RECT 1014.440 713.780 1015.560 717.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 674.580 1015.560 677.820 ;
  LAYER ME3 ;
  RECT 1014.440 674.580 1015.560 677.820 ;
  LAYER ME2 ;
  RECT 1014.440 674.580 1015.560 677.820 ;
  LAYER ME1 ;
  RECT 1014.440 674.580 1015.560 677.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 666.740 1015.560 669.980 ;
  LAYER ME3 ;
  RECT 1014.440 666.740 1015.560 669.980 ;
  LAYER ME2 ;
  RECT 1014.440 666.740 1015.560 669.980 ;
  LAYER ME1 ;
  RECT 1014.440 666.740 1015.560 669.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 658.900 1015.560 662.140 ;
  LAYER ME3 ;
  RECT 1014.440 658.900 1015.560 662.140 ;
  LAYER ME2 ;
  RECT 1014.440 658.900 1015.560 662.140 ;
  LAYER ME1 ;
  RECT 1014.440 658.900 1015.560 662.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 651.060 1015.560 654.300 ;
  LAYER ME3 ;
  RECT 1014.440 651.060 1015.560 654.300 ;
  LAYER ME2 ;
  RECT 1014.440 651.060 1015.560 654.300 ;
  LAYER ME1 ;
  RECT 1014.440 651.060 1015.560 654.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 643.220 1015.560 646.460 ;
  LAYER ME3 ;
  RECT 1014.440 643.220 1015.560 646.460 ;
  LAYER ME2 ;
  RECT 1014.440 643.220 1015.560 646.460 ;
  LAYER ME1 ;
  RECT 1014.440 643.220 1015.560 646.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 635.380 1015.560 638.620 ;
  LAYER ME3 ;
  RECT 1014.440 635.380 1015.560 638.620 ;
  LAYER ME2 ;
  RECT 1014.440 635.380 1015.560 638.620 ;
  LAYER ME1 ;
  RECT 1014.440 635.380 1015.560 638.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 596.180 1015.560 599.420 ;
  LAYER ME3 ;
  RECT 1014.440 596.180 1015.560 599.420 ;
  LAYER ME2 ;
  RECT 1014.440 596.180 1015.560 599.420 ;
  LAYER ME1 ;
  RECT 1014.440 596.180 1015.560 599.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 588.340 1015.560 591.580 ;
  LAYER ME3 ;
  RECT 1014.440 588.340 1015.560 591.580 ;
  LAYER ME2 ;
  RECT 1014.440 588.340 1015.560 591.580 ;
  LAYER ME1 ;
  RECT 1014.440 588.340 1015.560 591.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 580.500 1015.560 583.740 ;
  LAYER ME3 ;
  RECT 1014.440 580.500 1015.560 583.740 ;
  LAYER ME2 ;
  RECT 1014.440 580.500 1015.560 583.740 ;
  LAYER ME1 ;
  RECT 1014.440 580.500 1015.560 583.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 572.660 1015.560 575.900 ;
  LAYER ME3 ;
  RECT 1014.440 572.660 1015.560 575.900 ;
  LAYER ME2 ;
  RECT 1014.440 572.660 1015.560 575.900 ;
  LAYER ME1 ;
  RECT 1014.440 572.660 1015.560 575.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 564.820 1015.560 568.060 ;
  LAYER ME3 ;
  RECT 1014.440 564.820 1015.560 568.060 ;
  LAYER ME2 ;
  RECT 1014.440 564.820 1015.560 568.060 ;
  LAYER ME1 ;
  RECT 1014.440 564.820 1015.560 568.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 556.980 1015.560 560.220 ;
  LAYER ME3 ;
  RECT 1014.440 556.980 1015.560 560.220 ;
  LAYER ME2 ;
  RECT 1014.440 556.980 1015.560 560.220 ;
  LAYER ME1 ;
  RECT 1014.440 556.980 1015.560 560.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 517.780 1015.560 521.020 ;
  LAYER ME3 ;
  RECT 1014.440 517.780 1015.560 521.020 ;
  LAYER ME2 ;
  RECT 1014.440 517.780 1015.560 521.020 ;
  LAYER ME1 ;
  RECT 1014.440 517.780 1015.560 521.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 509.940 1015.560 513.180 ;
  LAYER ME3 ;
  RECT 1014.440 509.940 1015.560 513.180 ;
  LAYER ME2 ;
  RECT 1014.440 509.940 1015.560 513.180 ;
  LAYER ME1 ;
  RECT 1014.440 509.940 1015.560 513.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 502.100 1015.560 505.340 ;
  LAYER ME3 ;
  RECT 1014.440 502.100 1015.560 505.340 ;
  LAYER ME2 ;
  RECT 1014.440 502.100 1015.560 505.340 ;
  LAYER ME1 ;
  RECT 1014.440 502.100 1015.560 505.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 494.260 1015.560 497.500 ;
  LAYER ME3 ;
  RECT 1014.440 494.260 1015.560 497.500 ;
  LAYER ME2 ;
  RECT 1014.440 494.260 1015.560 497.500 ;
  LAYER ME1 ;
  RECT 1014.440 494.260 1015.560 497.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 486.420 1015.560 489.660 ;
  LAYER ME3 ;
  RECT 1014.440 486.420 1015.560 489.660 ;
  LAYER ME2 ;
  RECT 1014.440 486.420 1015.560 489.660 ;
  LAYER ME1 ;
  RECT 1014.440 486.420 1015.560 489.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 478.580 1015.560 481.820 ;
  LAYER ME3 ;
  RECT 1014.440 478.580 1015.560 481.820 ;
  LAYER ME2 ;
  RECT 1014.440 478.580 1015.560 481.820 ;
  LAYER ME1 ;
  RECT 1014.440 478.580 1015.560 481.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 439.380 1015.560 442.620 ;
  LAYER ME3 ;
  RECT 1014.440 439.380 1015.560 442.620 ;
  LAYER ME2 ;
  RECT 1014.440 439.380 1015.560 442.620 ;
  LAYER ME1 ;
  RECT 1014.440 439.380 1015.560 442.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 431.540 1015.560 434.780 ;
  LAYER ME3 ;
  RECT 1014.440 431.540 1015.560 434.780 ;
  LAYER ME2 ;
  RECT 1014.440 431.540 1015.560 434.780 ;
  LAYER ME1 ;
  RECT 1014.440 431.540 1015.560 434.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 423.700 1015.560 426.940 ;
  LAYER ME3 ;
  RECT 1014.440 423.700 1015.560 426.940 ;
  LAYER ME2 ;
  RECT 1014.440 423.700 1015.560 426.940 ;
  LAYER ME1 ;
  RECT 1014.440 423.700 1015.560 426.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 415.860 1015.560 419.100 ;
  LAYER ME3 ;
  RECT 1014.440 415.860 1015.560 419.100 ;
  LAYER ME2 ;
  RECT 1014.440 415.860 1015.560 419.100 ;
  LAYER ME1 ;
  RECT 1014.440 415.860 1015.560 419.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 408.020 1015.560 411.260 ;
  LAYER ME3 ;
  RECT 1014.440 408.020 1015.560 411.260 ;
  LAYER ME2 ;
  RECT 1014.440 408.020 1015.560 411.260 ;
  LAYER ME1 ;
  RECT 1014.440 408.020 1015.560 411.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 400.180 1015.560 403.420 ;
  LAYER ME3 ;
  RECT 1014.440 400.180 1015.560 403.420 ;
  LAYER ME2 ;
  RECT 1014.440 400.180 1015.560 403.420 ;
  LAYER ME1 ;
  RECT 1014.440 400.180 1015.560 403.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 360.980 1015.560 364.220 ;
  LAYER ME3 ;
  RECT 1014.440 360.980 1015.560 364.220 ;
  LAYER ME2 ;
  RECT 1014.440 360.980 1015.560 364.220 ;
  LAYER ME1 ;
  RECT 1014.440 360.980 1015.560 364.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 353.140 1015.560 356.380 ;
  LAYER ME3 ;
  RECT 1014.440 353.140 1015.560 356.380 ;
  LAYER ME2 ;
  RECT 1014.440 353.140 1015.560 356.380 ;
  LAYER ME1 ;
  RECT 1014.440 353.140 1015.560 356.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 345.300 1015.560 348.540 ;
  LAYER ME3 ;
  RECT 1014.440 345.300 1015.560 348.540 ;
  LAYER ME2 ;
  RECT 1014.440 345.300 1015.560 348.540 ;
  LAYER ME1 ;
  RECT 1014.440 345.300 1015.560 348.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 337.460 1015.560 340.700 ;
  LAYER ME3 ;
  RECT 1014.440 337.460 1015.560 340.700 ;
  LAYER ME2 ;
  RECT 1014.440 337.460 1015.560 340.700 ;
  LAYER ME1 ;
  RECT 1014.440 337.460 1015.560 340.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 329.620 1015.560 332.860 ;
  LAYER ME3 ;
  RECT 1014.440 329.620 1015.560 332.860 ;
  LAYER ME2 ;
  RECT 1014.440 329.620 1015.560 332.860 ;
  LAYER ME1 ;
  RECT 1014.440 329.620 1015.560 332.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 321.780 1015.560 325.020 ;
  LAYER ME3 ;
  RECT 1014.440 321.780 1015.560 325.020 ;
  LAYER ME2 ;
  RECT 1014.440 321.780 1015.560 325.020 ;
  LAYER ME1 ;
  RECT 1014.440 321.780 1015.560 325.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 282.580 1015.560 285.820 ;
  LAYER ME3 ;
  RECT 1014.440 282.580 1015.560 285.820 ;
  LAYER ME2 ;
  RECT 1014.440 282.580 1015.560 285.820 ;
  LAYER ME1 ;
  RECT 1014.440 282.580 1015.560 285.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 274.740 1015.560 277.980 ;
  LAYER ME3 ;
  RECT 1014.440 274.740 1015.560 277.980 ;
  LAYER ME2 ;
  RECT 1014.440 274.740 1015.560 277.980 ;
  LAYER ME1 ;
  RECT 1014.440 274.740 1015.560 277.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 266.900 1015.560 270.140 ;
  LAYER ME3 ;
  RECT 1014.440 266.900 1015.560 270.140 ;
  LAYER ME2 ;
  RECT 1014.440 266.900 1015.560 270.140 ;
  LAYER ME1 ;
  RECT 1014.440 266.900 1015.560 270.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 259.060 1015.560 262.300 ;
  LAYER ME3 ;
  RECT 1014.440 259.060 1015.560 262.300 ;
  LAYER ME2 ;
  RECT 1014.440 259.060 1015.560 262.300 ;
  LAYER ME1 ;
  RECT 1014.440 259.060 1015.560 262.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 251.220 1015.560 254.460 ;
  LAYER ME3 ;
  RECT 1014.440 251.220 1015.560 254.460 ;
  LAYER ME2 ;
  RECT 1014.440 251.220 1015.560 254.460 ;
  LAYER ME1 ;
  RECT 1014.440 251.220 1015.560 254.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 243.380 1015.560 246.620 ;
  LAYER ME3 ;
  RECT 1014.440 243.380 1015.560 246.620 ;
  LAYER ME2 ;
  RECT 1014.440 243.380 1015.560 246.620 ;
  LAYER ME1 ;
  RECT 1014.440 243.380 1015.560 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 204.180 1015.560 207.420 ;
  LAYER ME3 ;
  RECT 1014.440 204.180 1015.560 207.420 ;
  LAYER ME2 ;
  RECT 1014.440 204.180 1015.560 207.420 ;
  LAYER ME1 ;
  RECT 1014.440 204.180 1015.560 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 196.340 1015.560 199.580 ;
  LAYER ME3 ;
  RECT 1014.440 196.340 1015.560 199.580 ;
  LAYER ME2 ;
  RECT 1014.440 196.340 1015.560 199.580 ;
  LAYER ME1 ;
  RECT 1014.440 196.340 1015.560 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 188.500 1015.560 191.740 ;
  LAYER ME3 ;
  RECT 1014.440 188.500 1015.560 191.740 ;
  LAYER ME2 ;
  RECT 1014.440 188.500 1015.560 191.740 ;
  LAYER ME1 ;
  RECT 1014.440 188.500 1015.560 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 180.660 1015.560 183.900 ;
  LAYER ME3 ;
  RECT 1014.440 180.660 1015.560 183.900 ;
  LAYER ME2 ;
  RECT 1014.440 180.660 1015.560 183.900 ;
  LAYER ME1 ;
  RECT 1014.440 180.660 1015.560 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 172.820 1015.560 176.060 ;
  LAYER ME3 ;
  RECT 1014.440 172.820 1015.560 176.060 ;
  LAYER ME2 ;
  RECT 1014.440 172.820 1015.560 176.060 ;
  LAYER ME1 ;
  RECT 1014.440 172.820 1015.560 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 164.980 1015.560 168.220 ;
  LAYER ME3 ;
  RECT 1014.440 164.980 1015.560 168.220 ;
  LAYER ME2 ;
  RECT 1014.440 164.980 1015.560 168.220 ;
  LAYER ME1 ;
  RECT 1014.440 164.980 1015.560 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 125.780 1015.560 129.020 ;
  LAYER ME3 ;
  RECT 1014.440 125.780 1015.560 129.020 ;
  LAYER ME2 ;
  RECT 1014.440 125.780 1015.560 129.020 ;
  LAYER ME1 ;
  RECT 1014.440 125.780 1015.560 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 117.940 1015.560 121.180 ;
  LAYER ME3 ;
  RECT 1014.440 117.940 1015.560 121.180 ;
  LAYER ME2 ;
  RECT 1014.440 117.940 1015.560 121.180 ;
  LAYER ME1 ;
  RECT 1014.440 117.940 1015.560 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 110.100 1015.560 113.340 ;
  LAYER ME3 ;
  RECT 1014.440 110.100 1015.560 113.340 ;
  LAYER ME2 ;
  RECT 1014.440 110.100 1015.560 113.340 ;
  LAYER ME1 ;
  RECT 1014.440 110.100 1015.560 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 102.260 1015.560 105.500 ;
  LAYER ME3 ;
  RECT 1014.440 102.260 1015.560 105.500 ;
  LAYER ME2 ;
  RECT 1014.440 102.260 1015.560 105.500 ;
  LAYER ME1 ;
  RECT 1014.440 102.260 1015.560 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 94.420 1015.560 97.660 ;
  LAYER ME3 ;
  RECT 1014.440 94.420 1015.560 97.660 ;
  LAYER ME2 ;
  RECT 1014.440 94.420 1015.560 97.660 ;
  LAYER ME1 ;
  RECT 1014.440 94.420 1015.560 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 86.580 1015.560 89.820 ;
  LAYER ME3 ;
  RECT 1014.440 86.580 1015.560 89.820 ;
  LAYER ME2 ;
  RECT 1014.440 86.580 1015.560 89.820 ;
  LAYER ME1 ;
  RECT 1014.440 86.580 1015.560 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 47.380 1015.560 50.620 ;
  LAYER ME3 ;
  RECT 1014.440 47.380 1015.560 50.620 ;
  LAYER ME2 ;
  RECT 1014.440 47.380 1015.560 50.620 ;
  LAYER ME1 ;
  RECT 1014.440 47.380 1015.560 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 39.540 1015.560 42.780 ;
  LAYER ME3 ;
  RECT 1014.440 39.540 1015.560 42.780 ;
  LAYER ME2 ;
  RECT 1014.440 39.540 1015.560 42.780 ;
  LAYER ME1 ;
  RECT 1014.440 39.540 1015.560 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 31.700 1015.560 34.940 ;
  LAYER ME3 ;
  RECT 1014.440 31.700 1015.560 34.940 ;
  LAYER ME2 ;
  RECT 1014.440 31.700 1015.560 34.940 ;
  LAYER ME1 ;
  RECT 1014.440 31.700 1015.560 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 23.860 1015.560 27.100 ;
  LAYER ME3 ;
  RECT 1014.440 23.860 1015.560 27.100 ;
  LAYER ME2 ;
  RECT 1014.440 23.860 1015.560 27.100 ;
  LAYER ME1 ;
  RECT 1014.440 23.860 1015.560 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 16.020 1015.560 19.260 ;
  LAYER ME3 ;
  RECT 1014.440 16.020 1015.560 19.260 ;
  LAYER ME2 ;
  RECT 1014.440 16.020 1015.560 19.260 ;
  LAYER ME1 ;
  RECT 1014.440 16.020 1015.560 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 8.180 1015.560 11.420 ;
  LAYER ME3 ;
  RECT 1014.440 8.180 1015.560 11.420 ;
  LAYER ME2 ;
  RECT 1014.440 8.180 1015.560 11.420 ;
  LAYER ME1 ;
  RECT 1014.440 8.180 1015.560 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1380.180 1.120 1383.420 ;
  LAYER ME3 ;
  RECT 0.000 1380.180 1.120 1383.420 ;
  LAYER ME2 ;
  RECT 0.000 1380.180 1.120 1383.420 ;
  LAYER ME1 ;
  RECT 0.000 1380.180 1.120 1383.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1372.340 1.120 1375.580 ;
  LAYER ME3 ;
  RECT 0.000 1372.340 1.120 1375.580 ;
  LAYER ME2 ;
  RECT 0.000 1372.340 1.120 1375.580 ;
  LAYER ME1 ;
  RECT 0.000 1372.340 1.120 1375.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1364.500 1.120 1367.740 ;
  LAYER ME3 ;
  RECT 0.000 1364.500 1.120 1367.740 ;
  LAYER ME2 ;
  RECT 0.000 1364.500 1.120 1367.740 ;
  LAYER ME1 ;
  RECT 0.000 1364.500 1.120 1367.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1356.660 1.120 1359.900 ;
  LAYER ME3 ;
  RECT 0.000 1356.660 1.120 1359.900 ;
  LAYER ME2 ;
  RECT 0.000 1356.660 1.120 1359.900 ;
  LAYER ME1 ;
  RECT 0.000 1356.660 1.120 1359.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1348.820 1.120 1352.060 ;
  LAYER ME3 ;
  RECT 0.000 1348.820 1.120 1352.060 ;
  LAYER ME2 ;
  RECT 0.000 1348.820 1.120 1352.060 ;
  LAYER ME1 ;
  RECT 0.000 1348.820 1.120 1352.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1340.980 1.120 1344.220 ;
  LAYER ME3 ;
  RECT 0.000 1340.980 1.120 1344.220 ;
  LAYER ME2 ;
  RECT 0.000 1340.980 1.120 1344.220 ;
  LAYER ME1 ;
  RECT 0.000 1340.980 1.120 1344.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1301.780 1.120 1305.020 ;
  LAYER ME3 ;
  RECT 0.000 1301.780 1.120 1305.020 ;
  LAYER ME2 ;
  RECT 0.000 1301.780 1.120 1305.020 ;
  LAYER ME1 ;
  RECT 0.000 1301.780 1.120 1305.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1293.940 1.120 1297.180 ;
  LAYER ME3 ;
  RECT 0.000 1293.940 1.120 1297.180 ;
  LAYER ME2 ;
  RECT 0.000 1293.940 1.120 1297.180 ;
  LAYER ME1 ;
  RECT 0.000 1293.940 1.120 1297.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1286.100 1.120 1289.340 ;
  LAYER ME3 ;
  RECT 0.000 1286.100 1.120 1289.340 ;
  LAYER ME2 ;
  RECT 0.000 1286.100 1.120 1289.340 ;
  LAYER ME1 ;
  RECT 0.000 1286.100 1.120 1289.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1278.260 1.120 1281.500 ;
  LAYER ME3 ;
  RECT 0.000 1278.260 1.120 1281.500 ;
  LAYER ME2 ;
  RECT 0.000 1278.260 1.120 1281.500 ;
  LAYER ME1 ;
  RECT 0.000 1278.260 1.120 1281.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1270.420 1.120 1273.660 ;
  LAYER ME3 ;
  RECT 0.000 1270.420 1.120 1273.660 ;
  LAYER ME2 ;
  RECT 0.000 1270.420 1.120 1273.660 ;
  LAYER ME1 ;
  RECT 0.000 1270.420 1.120 1273.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1262.580 1.120 1265.820 ;
  LAYER ME3 ;
  RECT 0.000 1262.580 1.120 1265.820 ;
  LAYER ME2 ;
  RECT 0.000 1262.580 1.120 1265.820 ;
  LAYER ME1 ;
  RECT 0.000 1262.580 1.120 1265.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1223.380 1.120 1226.620 ;
  LAYER ME3 ;
  RECT 0.000 1223.380 1.120 1226.620 ;
  LAYER ME2 ;
  RECT 0.000 1223.380 1.120 1226.620 ;
  LAYER ME1 ;
  RECT 0.000 1223.380 1.120 1226.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1215.540 1.120 1218.780 ;
  LAYER ME3 ;
  RECT 0.000 1215.540 1.120 1218.780 ;
  LAYER ME2 ;
  RECT 0.000 1215.540 1.120 1218.780 ;
  LAYER ME1 ;
  RECT 0.000 1215.540 1.120 1218.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1207.700 1.120 1210.940 ;
  LAYER ME3 ;
  RECT 0.000 1207.700 1.120 1210.940 ;
  LAYER ME2 ;
  RECT 0.000 1207.700 1.120 1210.940 ;
  LAYER ME1 ;
  RECT 0.000 1207.700 1.120 1210.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1199.860 1.120 1203.100 ;
  LAYER ME3 ;
  RECT 0.000 1199.860 1.120 1203.100 ;
  LAYER ME2 ;
  RECT 0.000 1199.860 1.120 1203.100 ;
  LAYER ME1 ;
  RECT 0.000 1199.860 1.120 1203.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1192.020 1.120 1195.260 ;
  LAYER ME3 ;
  RECT 0.000 1192.020 1.120 1195.260 ;
  LAYER ME2 ;
  RECT 0.000 1192.020 1.120 1195.260 ;
  LAYER ME1 ;
  RECT 0.000 1192.020 1.120 1195.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1184.180 1.120 1187.420 ;
  LAYER ME3 ;
  RECT 0.000 1184.180 1.120 1187.420 ;
  LAYER ME2 ;
  RECT 0.000 1184.180 1.120 1187.420 ;
  LAYER ME1 ;
  RECT 0.000 1184.180 1.120 1187.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1144.980 1.120 1148.220 ;
  LAYER ME3 ;
  RECT 0.000 1144.980 1.120 1148.220 ;
  LAYER ME2 ;
  RECT 0.000 1144.980 1.120 1148.220 ;
  LAYER ME1 ;
  RECT 0.000 1144.980 1.120 1148.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1137.140 1.120 1140.380 ;
  LAYER ME3 ;
  RECT 0.000 1137.140 1.120 1140.380 ;
  LAYER ME2 ;
  RECT 0.000 1137.140 1.120 1140.380 ;
  LAYER ME1 ;
  RECT 0.000 1137.140 1.120 1140.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1129.300 1.120 1132.540 ;
  LAYER ME3 ;
  RECT 0.000 1129.300 1.120 1132.540 ;
  LAYER ME2 ;
  RECT 0.000 1129.300 1.120 1132.540 ;
  LAYER ME1 ;
  RECT 0.000 1129.300 1.120 1132.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1121.460 1.120 1124.700 ;
  LAYER ME3 ;
  RECT 0.000 1121.460 1.120 1124.700 ;
  LAYER ME2 ;
  RECT 0.000 1121.460 1.120 1124.700 ;
  LAYER ME1 ;
  RECT 0.000 1121.460 1.120 1124.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1113.620 1.120 1116.860 ;
  LAYER ME3 ;
  RECT 0.000 1113.620 1.120 1116.860 ;
  LAYER ME2 ;
  RECT 0.000 1113.620 1.120 1116.860 ;
  LAYER ME1 ;
  RECT 0.000 1113.620 1.120 1116.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1105.780 1.120 1109.020 ;
  LAYER ME3 ;
  RECT 0.000 1105.780 1.120 1109.020 ;
  LAYER ME2 ;
  RECT 0.000 1105.780 1.120 1109.020 ;
  LAYER ME1 ;
  RECT 0.000 1105.780 1.120 1109.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER ME3 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER ME2 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER ME1 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER ME3 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER ME2 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER ME1 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER ME3 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER ME2 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER ME1 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER ME3 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER ME2 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER ME1 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER ME3 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER ME2 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER ME1 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER ME3 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER ME2 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER ME1 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER ME3 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER ME2 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER ME1 ;
  RECT 0.000 988.180 1.120 991.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER ME3 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER ME2 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER ME1 ;
  RECT 0.000 980.340 1.120 983.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER ME3 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER ME2 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER ME1 ;
  RECT 0.000 972.500 1.120 975.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER ME3 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER ME2 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER ME1 ;
  RECT 0.000 964.660 1.120 967.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER ME3 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER ME2 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER ME1 ;
  RECT 0.000 956.820 1.120 960.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER ME3 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER ME2 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER ME1 ;
  RECT 0.000 948.980 1.120 952.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER ME3 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER ME2 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER ME1 ;
  RECT 0.000 909.780 1.120 913.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER ME3 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER ME2 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER ME1 ;
  RECT 0.000 901.940 1.120 905.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER ME3 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER ME2 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER ME1 ;
  RECT 0.000 894.100 1.120 897.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER ME3 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER ME2 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER ME1 ;
  RECT 0.000 886.260 1.120 889.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER ME3 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER ME2 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER ME1 ;
  RECT 0.000 878.420 1.120 881.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER ME3 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER ME2 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER ME1 ;
  RECT 0.000 870.580 1.120 873.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER ME3 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER ME2 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER ME1 ;
  RECT 0.000 831.380 1.120 834.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER ME3 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER ME2 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER ME1 ;
  RECT 0.000 823.540 1.120 826.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER ME3 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER ME2 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER ME1 ;
  RECT 0.000 815.700 1.120 818.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER ME3 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER ME2 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER ME1 ;
  RECT 0.000 807.860 1.120 811.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER ME3 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER ME2 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER ME1 ;
  RECT 0.000 800.020 1.120 803.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER ME3 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER ME2 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER ME1 ;
  RECT 0.000 792.180 1.120 795.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER ME3 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER ME2 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER ME1 ;
  RECT 0.000 752.980 1.120 756.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER ME3 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER ME2 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER ME1 ;
  RECT 0.000 745.140 1.120 748.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER ME3 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER ME2 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER ME1 ;
  RECT 0.000 737.300 1.120 740.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER ME3 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER ME2 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER ME1 ;
  RECT 0.000 729.460 1.120 732.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER ME3 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER ME2 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER ME1 ;
  RECT 0.000 721.620 1.120 724.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER ME3 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER ME2 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER ME1 ;
  RECT 0.000 713.780 1.120 717.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER ME3 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER ME2 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER ME1 ;
  RECT 0.000 674.580 1.120 677.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER ME3 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER ME2 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER ME1 ;
  RECT 0.000 666.740 1.120 669.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER ME3 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER ME2 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER ME1 ;
  RECT 0.000 658.900 1.120 662.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER ME3 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER ME2 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER ME1 ;
  RECT 0.000 651.060 1.120 654.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER ME3 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER ME2 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER ME1 ;
  RECT 0.000 643.220 1.120 646.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER ME3 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER ME2 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER ME1 ;
  RECT 0.000 635.380 1.120 638.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER ME3 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER ME2 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER ME1 ;
  RECT 0.000 596.180 1.120 599.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER ME3 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER ME2 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER ME1 ;
  RECT 0.000 588.340 1.120 591.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER ME3 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER ME2 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER ME1 ;
  RECT 0.000 580.500 1.120 583.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER ME3 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER ME2 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER ME1 ;
  RECT 0.000 572.660 1.120 575.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER ME3 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER ME2 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER ME1 ;
  RECT 0.000 564.820 1.120 568.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER ME3 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER ME2 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER ME1 ;
  RECT 0.000 556.980 1.120 560.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER ME3 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER ME2 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER ME1 ;
  RECT 0.000 517.780 1.120 521.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER ME3 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER ME2 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER ME1 ;
  RECT 0.000 509.940 1.120 513.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER ME3 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER ME2 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER ME1 ;
  RECT 0.000 502.100 1.120 505.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER ME3 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER ME2 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER ME1 ;
  RECT 0.000 494.260 1.120 497.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER ME3 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER ME2 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER ME1 ;
  RECT 0.000 486.420 1.120 489.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER ME3 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER ME2 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER ME1 ;
  RECT 0.000 478.580 1.120 481.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER ME3 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER ME2 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER ME1 ;
  RECT 0.000 439.380 1.120 442.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER ME3 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER ME2 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER ME1 ;
  RECT 0.000 431.540 1.120 434.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER ME3 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER ME2 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER ME1 ;
  RECT 0.000 423.700 1.120 426.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER ME3 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER ME2 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER ME1 ;
  RECT 0.000 415.860 1.120 419.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER ME3 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER ME2 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER ME1 ;
  RECT 0.000 408.020 1.120 411.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER ME3 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER ME2 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER ME1 ;
  RECT 0.000 400.180 1.120 403.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER ME3 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER ME2 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER ME1 ;
  RECT 0.000 360.980 1.120 364.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER ME3 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER ME2 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER ME1 ;
  RECT 0.000 353.140 1.120 356.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER ME3 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER ME2 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER ME1 ;
  RECT 0.000 345.300 1.120 348.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER ME3 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER ME2 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER ME1 ;
  RECT 0.000 337.460 1.120 340.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER ME3 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER ME2 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER ME1 ;
  RECT 0.000 329.620 1.120 332.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER ME3 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER ME2 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER ME1 ;
  RECT 0.000 321.780 1.120 325.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 997.360 1390.480 1000.900 1391.600 ;
  LAYER ME3 ;
  RECT 997.360 1390.480 1000.900 1391.600 ;
  LAYER ME2 ;
  RECT 997.360 1390.480 1000.900 1391.600 ;
  LAYER ME1 ;
  RECT 997.360 1390.480 1000.900 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 988.680 1390.480 992.220 1391.600 ;
  LAYER ME3 ;
  RECT 988.680 1390.480 992.220 1391.600 ;
  LAYER ME2 ;
  RECT 988.680 1390.480 992.220 1391.600 ;
  LAYER ME1 ;
  RECT 988.680 1390.480 992.220 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 980.000 1390.480 983.540 1391.600 ;
  LAYER ME3 ;
  RECT 980.000 1390.480 983.540 1391.600 ;
  LAYER ME2 ;
  RECT 980.000 1390.480 983.540 1391.600 ;
  LAYER ME1 ;
  RECT 980.000 1390.480 983.540 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 971.320 1390.480 974.860 1391.600 ;
  LAYER ME3 ;
  RECT 971.320 1390.480 974.860 1391.600 ;
  LAYER ME2 ;
  RECT 971.320 1390.480 974.860 1391.600 ;
  LAYER ME1 ;
  RECT 971.320 1390.480 974.860 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 962.640 1390.480 966.180 1391.600 ;
  LAYER ME3 ;
  RECT 962.640 1390.480 966.180 1391.600 ;
  LAYER ME2 ;
  RECT 962.640 1390.480 966.180 1391.600 ;
  LAYER ME1 ;
  RECT 962.640 1390.480 966.180 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 919.240 1390.480 922.780 1391.600 ;
  LAYER ME3 ;
  RECT 919.240 1390.480 922.780 1391.600 ;
  LAYER ME2 ;
  RECT 919.240 1390.480 922.780 1391.600 ;
  LAYER ME1 ;
  RECT 919.240 1390.480 922.780 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 910.560 1390.480 914.100 1391.600 ;
  LAYER ME3 ;
  RECT 910.560 1390.480 914.100 1391.600 ;
  LAYER ME2 ;
  RECT 910.560 1390.480 914.100 1391.600 ;
  LAYER ME1 ;
  RECT 910.560 1390.480 914.100 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 901.880 1390.480 905.420 1391.600 ;
  LAYER ME3 ;
  RECT 901.880 1390.480 905.420 1391.600 ;
  LAYER ME2 ;
  RECT 901.880 1390.480 905.420 1391.600 ;
  LAYER ME1 ;
  RECT 901.880 1390.480 905.420 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 893.200 1390.480 896.740 1391.600 ;
  LAYER ME3 ;
  RECT 893.200 1390.480 896.740 1391.600 ;
  LAYER ME2 ;
  RECT 893.200 1390.480 896.740 1391.600 ;
  LAYER ME1 ;
  RECT 893.200 1390.480 896.740 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 884.520 1390.480 888.060 1391.600 ;
  LAYER ME3 ;
  RECT 884.520 1390.480 888.060 1391.600 ;
  LAYER ME2 ;
  RECT 884.520 1390.480 888.060 1391.600 ;
  LAYER ME1 ;
  RECT 884.520 1390.480 888.060 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 875.840 1390.480 879.380 1391.600 ;
  LAYER ME3 ;
  RECT 875.840 1390.480 879.380 1391.600 ;
  LAYER ME2 ;
  RECT 875.840 1390.480 879.380 1391.600 ;
  LAYER ME1 ;
  RECT 875.840 1390.480 879.380 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 832.440 1390.480 835.980 1391.600 ;
  LAYER ME3 ;
  RECT 832.440 1390.480 835.980 1391.600 ;
  LAYER ME2 ;
  RECT 832.440 1390.480 835.980 1391.600 ;
  LAYER ME1 ;
  RECT 832.440 1390.480 835.980 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 823.760 1390.480 827.300 1391.600 ;
  LAYER ME3 ;
  RECT 823.760 1390.480 827.300 1391.600 ;
  LAYER ME2 ;
  RECT 823.760 1390.480 827.300 1391.600 ;
  LAYER ME1 ;
  RECT 823.760 1390.480 827.300 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 815.080 1390.480 818.620 1391.600 ;
  LAYER ME3 ;
  RECT 815.080 1390.480 818.620 1391.600 ;
  LAYER ME2 ;
  RECT 815.080 1390.480 818.620 1391.600 ;
  LAYER ME1 ;
  RECT 815.080 1390.480 818.620 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 806.400 1390.480 809.940 1391.600 ;
  LAYER ME3 ;
  RECT 806.400 1390.480 809.940 1391.600 ;
  LAYER ME2 ;
  RECT 806.400 1390.480 809.940 1391.600 ;
  LAYER ME1 ;
  RECT 806.400 1390.480 809.940 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 797.720 1390.480 801.260 1391.600 ;
  LAYER ME3 ;
  RECT 797.720 1390.480 801.260 1391.600 ;
  LAYER ME2 ;
  RECT 797.720 1390.480 801.260 1391.600 ;
  LAYER ME1 ;
  RECT 797.720 1390.480 801.260 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 789.040 1390.480 792.580 1391.600 ;
  LAYER ME3 ;
  RECT 789.040 1390.480 792.580 1391.600 ;
  LAYER ME2 ;
  RECT 789.040 1390.480 792.580 1391.600 ;
  LAYER ME1 ;
  RECT 789.040 1390.480 792.580 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 745.640 1390.480 749.180 1391.600 ;
  LAYER ME3 ;
  RECT 745.640 1390.480 749.180 1391.600 ;
  LAYER ME2 ;
  RECT 745.640 1390.480 749.180 1391.600 ;
  LAYER ME1 ;
  RECT 745.640 1390.480 749.180 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 736.960 1390.480 740.500 1391.600 ;
  LAYER ME3 ;
  RECT 736.960 1390.480 740.500 1391.600 ;
  LAYER ME2 ;
  RECT 736.960 1390.480 740.500 1391.600 ;
  LAYER ME1 ;
  RECT 736.960 1390.480 740.500 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 728.280 1390.480 731.820 1391.600 ;
  LAYER ME3 ;
  RECT 728.280 1390.480 731.820 1391.600 ;
  LAYER ME2 ;
  RECT 728.280 1390.480 731.820 1391.600 ;
  LAYER ME1 ;
  RECT 728.280 1390.480 731.820 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 719.600 1390.480 723.140 1391.600 ;
  LAYER ME3 ;
  RECT 719.600 1390.480 723.140 1391.600 ;
  LAYER ME2 ;
  RECT 719.600 1390.480 723.140 1391.600 ;
  LAYER ME1 ;
  RECT 719.600 1390.480 723.140 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 710.920 1390.480 714.460 1391.600 ;
  LAYER ME3 ;
  RECT 710.920 1390.480 714.460 1391.600 ;
  LAYER ME2 ;
  RECT 710.920 1390.480 714.460 1391.600 ;
  LAYER ME1 ;
  RECT 710.920 1390.480 714.460 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 702.240 1390.480 705.780 1391.600 ;
  LAYER ME3 ;
  RECT 702.240 1390.480 705.780 1391.600 ;
  LAYER ME2 ;
  RECT 702.240 1390.480 705.780 1391.600 ;
  LAYER ME1 ;
  RECT 702.240 1390.480 705.780 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 658.840 1390.480 662.380 1391.600 ;
  LAYER ME3 ;
  RECT 658.840 1390.480 662.380 1391.600 ;
  LAYER ME2 ;
  RECT 658.840 1390.480 662.380 1391.600 ;
  LAYER ME1 ;
  RECT 658.840 1390.480 662.380 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 650.160 1390.480 653.700 1391.600 ;
  LAYER ME3 ;
  RECT 650.160 1390.480 653.700 1391.600 ;
  LAYER ME2 ;
  RECT 650.160 1390.480 653.700 1391.600 ;
  LAYER ME1 ;
  RECT 650.160 1390.480 653.700 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 641.480 1390.480 645.020 1391.600 ;
  LAYER ME3 ;
  RECT 641.480 1390.480 645.020 1391.600 ;
  LAYER ME2 ;
  RECT 641.480 1390.480 645.020 1391.600 ;
  LAYER ME1 ;
  RECT 641.480 1390.480 645.020 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 632.800 1390.480 636.340 1391.600 ;
  LAYER ME3 ;
  RECT 632.800 1390.480 636.340 1391.600 ;
  LAYER ME2 ;
  RECT 632.800 1390.480 636.340 1391.600 ;
  LAYER ME1 ;
  RECT 632.800 1390.480 636.340 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 624.120 1390.480 627.660 1391.600 ;
  LAYER ME3 ;
  RECT 624.120 1390.480 627.660 1391.600 ;
  LAYER ME2 ;
  RECT 624.120 1390.480 627.660 1391.600 ;
  LAYER ME1 ;
  RECT 624.120 1390.480 627.660 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 615.440 1390.480 618.980 1391.600 ;
  LAYER ME3 ;
  RECT 615.440 1390.480 618.980 1391.600 ;
  LAYER ME2 ;
  RECT 615.440 1390.480 618.980 1391.600 ;
  LAYER ME1 ;
  RECT 615.440 1390.480 618.980 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 572.040 1390.480 575.580 1391.600 ;
  LAYER ME3 ;
  RECT 572.040 1390.480 575.580 1391.600 ;
  LAYER ME2 ;
  RECT 572.040 1390.480 575.580 1391.600 ;
  LAYER ME1 ;
  RECT 572.040 1390.480 575.580 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 563.360 1390.480 566.900 1391.600 ;
  LAYER ME3 ;
  RECT 563.360 1390.480 566.900 1391.600 ;
  LAYER ME2 ;
  RECT 563.360 1390.480 566.900 1391.600 ;
  LAYER ME1 ;
  RECT 563.360 1390.480 566.900 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 554.680 1390.480 558.220 1391.600 ;
  LAYER ME3 ;
  RECT 554.680 1390.480 558.220 1391.600 ;
  LAYER ME2 ;
  RECT 554.680 1390.480 558.220 1391.600 ;
  LAYER ME1 ;
  RECT 554.680 1390.480 558.220 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.000 1390.480 549.540 1391.600 ;
  LAYER ME3 ;
  RECT 546.000 1390.480 549.540 1391.600 ;
  LAYER ME2 ;
  RECT 546.000 1390.480 549.540 1391.600 ;
  LAYER ME1 ;
  RECT 546.000 1390.480 549.540 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.320 1390.480 540.860 1391.600 ;
  LAYER ME3 ;
  RECT 537.320 1390.480 540.860 1391.600 ;
  LAYER ME2 ;
  RECT 537.320 1390.480 540.860 1391.600 ;
  LAYER ME1 ;
  RECT 537.320 1390.480 540.860 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.640 1390.480 532.180 1391.600 ;
  LAYER ME3 ;
  RECT 528.640 1390.480 532.180 1391.600 ;
  LAYER ME2 ;
  RECT 528.640 1390.480 532.180 1391.600 ;
  LAYER ME1 ;
  RECT 528.640 1390.480 532.180 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.240 1390.480 488.780 1391.600 ;
  LAYER ME3 ;
  RECT 485.240 1390.480 488.780 1391.600 ;
  LAYER ME2 ;
  RECT 485.240 1390.480 488.780 1391.600 ;
  LAYER ME1 ;
  RECT 485.240 1390.480 488.780 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.560 1390.480 480.100 1391.600 ;
  LAYER ME3 ;
  RECT 476.560 1390.480 480.100 1391.600 ;
  LAYER ME2 ;
  RECT 476.560 1390.480 480.100 1391.600 ;
  LAYER ME1 ;
  RECT 476.560 1390.480 480.100 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.880 1390.480 471.420 1391.600 ;
  LAYER ME3 ;
  RECT 467.880 1390.480 471.420 1391.600 ;
  LAYER ME2 ;
  RECT 467.880 1390.480 471.420 1391.600 ;
  LAYER ME1 ;
  RECT 467.880 1390.480 471.420 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.200 1390.480 462.740 1391.600 ;
  LAYER ME3 ;
  RECT 459.200 1390.480 462.740 1391.600 ;
  LAYER ME2 ;
  RECT 459.200 1390.480 462.740 1391.600 ;
  LAYER ME1 ;
  RECT 459.200 1390.480 462.740 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.520 1390.480 454.060 1391.600 ;
  LAYER ME3 ;
  RECT 450.520 1390.480 454.060 1391.600 ;
  LAYER ME2 ;
  RECT 450.520 1390.480 454.060 1391.600 ;
  LAYER ME1 ;
  RECT 450.520 1390.480 454.060 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.840 1390.480 445.380 1391.600 ;
  LAYER ME3 ;
  RECT 441.840 1390.480 445.380 1391.600 ;
  LAYER ME2 ;
  RECT 441.840 1390.480 445.380 1391.600 ;
  LAYER ME1 ;
  RECT 441.840 1390.480 445.380 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.440 1390.480 401.980 1391.600 ;
  LAYER ME3 ;
  RECT 398.440 1390.480 401.980 1391.600 ;
  LAYER ME2 ;
  RECT 398.440 1390.480 401.980 1391.600 ;
  LAYER ME1 ;
  RECT 398.440 1390.480 401.980 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.760 1390.480 393.300 1391.600 ;
  LAYER ME3 ;
  RECT 389.760 1390.480 393.300 1391.600 ;
  LAYER ME2 ;
  RECT 389.760 1390.480 393.300 1391.600 ;
  LAYER ME1 ;
  RECT 389.760 1390.480 393.300 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.080 1390.480 384.620 1391.600 ;
  LAYER ME3 ;
  RECT 381.080 1390.480 384.620 1391.600 ;
  LAYER ME2 ;
  RECT 381.080 1390.480 384.620 1391.600 ;
  LAYER ME1 ;
  RECT 381.080 1390.480 384.620 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.400 1390.480 375.940 1391.600 ;
  LAYER ME3 ;
  RECT 372.400 1390.480 375.940 1391.600 ;
  LAYER ME2 ;
  RECT 372.400 1390.480 375.940 1391.600 ;
  LAYER ME1 ;
  RECT 372.400 1390.480 375.940 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 1390.480 367.260 1391.600 ;
  LAYER ME3 ;
  RECT 363.720 1390.480 367.260 1391.600 ;
  LAYER ME2 ;
  RECT 363.720 1390.480 367.260 1391.600 ;
  LAYER ME1 ;
  RECT 363.720 1390.480 367.260 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.040 1390.480 358.580 1391.600 ;
  LAYER ME3 ;
  RECT 355.040 1390.480 358.580 1391.600 ;
  LAYER ME2 ;
  RECT 355.040 1390.480 358.580 1391.600 ;
  LAYER ME1 ;
  RECT 355.040 1390.480 358.580 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 1390.480 315.180 1391.600 ;
  LAYER ME3 ;
  RECT 311.640 1390.480 315.180 1391.600 ;
  LAYER ME2 ;
  RECT 311.640 1390.480 315.180 1391.600 ;
  LAYER ME1 ;
  RECT 311.640 1390.480 315.180 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 1390.480 306.500 1391.600 ;
  LAYER ME3 ;
  RECT 302.960 1390.480 306.500 1391.600 ;
  LAYER ME2 ;
  RECT 302.960 1390.480 306.500 1391.600 ;
  LAYER ME1 ;
  RECT 302.960 1390.480 306.500 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 1390.480 297.820 1391.600 ;
  LAYER ME3 ;
  RECT 294.280 1390.480 297.820 1391.600 ;
  LAYER ME2 ;
  RECT 294.280 1390.480 297.820 1391.600 ;
  LAYER ME1 ;
  RECT 294.280 1390.480 297.820 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 1390.480 289.140 1391.600 ;
  LAYER ME3 ;
  RECT 285.600 1390.480 289.140 1391.600 ;
  LAYER ME2 ;
  RECT 285.600 1390.480 289.140 1391.600 ;
  LAYER ME1 ;
  RECT 285.600 1390.480 289.140 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 1390.480 280.460 1391.600 ;
  LAYER ME3 ;
  RECT 276.920 1390.480 280.460 1391.600 ;
  LAYER ME2 ;
  RECT 276.920 1390.480 280.460 1391.600 ;
  LAYER ME1 ;
  RECT 276.920 1390.480 280.460 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 1390.480 271.780 1391.600 ;
  LAYER ME3 ;
  RECT 268.240 1390.480 271.780 1391.600 ;
  LAYER ME2 ;
  RECT 268.240 1390.480 271.780 1391.600 ;
  LAYER ME1 ;
  RECT 268.240 1390.480 271.780 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 1390.480 228.380 1391.600 ;
  LAYER ME3 ;
  RECT 224.840 1390.480 228.380 1391.600 ;
  LAYER ME2 ;
  RECT 224.840 1390.480 228.380 1391.600 ;
  LAYER ME1 ;
  RECT 224.840 1390.480 228.380 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 1390.480 219.700 1391.600 ;
  LAYER ME3 ;
  RECT 216.160 1390.480 219.700 1391.600 ;
  LAYER ME2 ;
  RECT 216.160 1390.480 219.700 1391.600 ;
  LAYER ME1 ;
  RECT 216.160 1390.480 219.700 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 1390.480 211.020 1391.600 ;
  LAYER ME3 ;
  RECT 207.480 1390.480 211.020 1391.600 ;
  LAYER ME2 ;
  RECT 207.480 1390.480 211.020 1391.600 ;
  LAYER ME1 ;
  RECT 207.480 1390.480 211.020 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 1390.480 202.340 1391.600 ;
  LAYER ME3 ;
  RECT 198.800 1390.480 202.340 1391.600 ;
  LAYER ME2 ;
  RECT 198.800 1390.480 202.340 1391.600 ;
  LAYER ME1 ;
  RECT 198.800 1390.480 202.340 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 1390.480 193.660 1391.600 ;
  LAYER ME3 ;
  RECT 190.120 1390.480 193.660 1391.600 ;
  LAYER ME2 ;
  RECT 190.120 1390.480 193.660 1391.600 ;
  LAYER ME1 ;
  RECT 190.120 1390.480 193.660 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 1390.480 184.980 1391.600 ;
  LAYER ME3 ;
  RECT 181.440 1390.480 184.980 1391.600 ;
  LAYER ME2 ;
  RECT 181.440 1390.480 184.980 1391.600 ;
  LAYER ME1 ;
  RECT 181.440 1390.480 184.980 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 1390.480 141.580 1391.600 ;
  LAYER ME3 ;
  RECT 138.040 1390.480 141.580 1391.600 ;
  LAYER ME2 ;
  RECT 138.040 1390.480 141.580 1391.600 ;
  LAYER ME1 ;
  RECT 138.040 1390.480 141.580 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 1390.480 132.900 1391.600 ;
  LAYER ME3 ;
  RECT 129.360 1390.480 132.900 1391.600 ;
  LAYER ME2 ;
  RECT 129.360 1390.480 132.900 1391.600 ;
  LAYER ME1 ;
  RECT 129.360 1390.480 132.900 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 1390.480 124.220 1391.600 ;
  LAYER ME3 ;
  RECT 120.680 1390.480 124.220 1391.600 ;
  LAYER ME2 ;
  RECT 120.680 1390.480 124.220 1391.600 ;
  LAYER ME1 ;
  RECT 120.680 1390.480 124.220 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 1390.480 115.540 1391.600 ;
  LAYER ME3 ;
  RECT 112.000 1390.480 115.540 1391.600 ;
  LAYER ME2 ;
  RECT 112.000 1390.480 115.540 1391.600 ;
  LAYER ME1 ;
  RECT 112.000 1390.480 115.540 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 1390.480 106.860 1391.600 ;
  LAYER ME3 ;
  RECT 103.320 1390.480 106.860 1391.600 ;
  LAYER ME2 ;
  RECT 103.320 1390.480 106.860 1391.600 ;
  LAYER ME1 ;
  RECT 103.320 1390.480 106.860 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 1390.480 98.180 1391.600 ;
  LAYER ME3 ;
  RECT 94.640 1390.480 98.180 1391.600 ;
  LAYER ME2 ;
  RECT 94.640 1390.480 98.180 1391.600 ;
  LAYER ME1 ;
  RECT 94.640 1390.480 98.180 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 1390.480 54.780 1391.600 ;
  LAYER ME3 ;
  RECT 51.240 1390.480 54.780 1391.600 ;
  LAYER ME2 ;
  RECT 51.240 1390.480 54.780 1391.600 ;
  LAYER ME1 ;
  RECT 51.240 1390.480 54.780 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 1390.480 46.100 1391.600 ;
  LAYER ME3 ;
  RECT 42.560 1390.480 46.100 1391.600 ;
  LAYER ME2 ;
  RECT 42.560 1390.480 46.100 1391.600 ;
  LAYER ME1 ;
  RECT 42.560 1390.480 46.100 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 1390.480 37.420 1391.600 ;
  LAYER ME3 ;
  RECT 33.880 1390.480 37.420 1391.600 ;
  LAYER ME2 ;
  RECT 33.880 1390.480 37.420 1391.600 ;
  LAYER ME1 ;
  RECT 33.880 1390.480 37.420 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 1390.480 28.740 1391.600 ;
  LAYER ME3 ;
  RECT 25.200 1390.480 28.740 1391.600 ;
  LAYER ME2 ;
  RECT 25.200 1390.480 28.740 1391.600 ;
  LAYER ME1 ;
  RECT 25.200 1390.480 28.740 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 1390.480 20.060 1391.600 ;
  LAYER ME3 ;
  RECT 16.520 1390.480 20.060 1391.600 ;
  LAYER ME2 ;
  RECT 16.520 1390.480 20.060 1391.600 ;
  LAYER ME1 ;
  RECT 16.520 1390.480 20.060 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 1390.480 11.380 1391.600 ;
  LAYER ME3 ;
  RECT 7.840 1390.480 11.380 1391.600 ;
  LAYER ME2 ;
  RECT 7.840 1390.480 11.380 1391.600 ;
  LAYER ME1 ;
  RECT 7.840 1390.480 11.380 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER ME3 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER ME2 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER ME1 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 991.780 0.000 995.320 1.120 ;
  LAYER ME3 ;
  RECT 991.780 0.000 995.320 1.120 ;
  LAYER ME2 ;
  RECT 991.780 0.000 995.320 1.120 ;
  LAYER ME1 ;
  RECT 991.780 0.000 995.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 983.100 0.000 986.640 1.120 ;
  LAYER ME3 ;
  RECT 983.100 0.000 986.640 1.120 ;
  LAYER ME2 ;
  RECT 983.100 0.000 986.640 1.120 ;
  LAYER ME1 ;
  RECT 983.100 0.000 986.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 974.420 0.000 977.960 1.120 ;
  LAYER ME3 ;
  RECT 974.420 0.000 977.960 1.120 ;
  LAYER ME2 ;
  RECT 974.420 0.000 977.960 1.120 ;
  LAYER ME1 ;
  RECT 974.420 0.000 977.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 952.720 0.000 956.260 1.120 ;
  LAYER ME3 ;
  RECT 952.720 0.000 956.260 1.120 ;
  LAYER ME2 ;
  RECT 952.720 0.000 956.260 1.120 ;
  LAYER ME1 ;
  RECT 952.720 0.000 956.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER ME3 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER ME2 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER ME1 ;
  RECT 887.620 0.000 891.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER ME3 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER ME2 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER ME1 ;
  RECT 878.940 0.000 882.480 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER ME3 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER ME2 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER ME1 ;
  RECT 870.260 0.000 873.800 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER ME3 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER ME2 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER ME1 ;
  RECT 861.580 0.000 865.120 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 839.880 0.000 843.420 1.120 ;
  LAYER ME3 ;
  RECT 839.880 0.000 843.420 1.120 ;
  LAYER ME2 ;
  RECT 839.880 0.000 843.420 1.120 ;
  LAYER ME1 ;
  RECT 839.880 0.000 843.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 826.240 0.000 829.780 1.120 ;
  LAYER ME3 ;
  RECT 826.240 0.000 829.780 1.120 ;
  LAYER ME2 ;
  RECT 826.240 0.000 829.780 1.120 ;
  LAYER ME1 ;
  RECT 826.240 0.000 829.780 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER ME3 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER ME2 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER ME1 ;
  RECT 761.140 0.000 764.680 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER ME3 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER ME2 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER ME1 ;
  RECT 752.460 0.000 756.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER ME3 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER ME2 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER ME1 ;
  RECT 740.060 0.000 743.600 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 717.740 0.000 721.280 1.120 ;
  LAYER ME3 ;
  RECT 717.740 0.000 721.280 1.120 ;
  LAYER ME2 ;
  RECT 717.740 0.000 721.280 1.120 ;
  LAYER ME1 ;
  RECT 717.740 0.000 721.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 709.060 0.000 712.600 1.120 ;
  LAYER ME3 ;
  RECT 709.060 0.000 712.600 1.120 ;
  LAYER ME2 ;
  RECT 709.060 0.000 712.600 1.120 ;
  LAYER ME1 ;
  RECT 709.060 0.000 712.600 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER ME3 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER ME2 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER ME1 ;
  RECT 700.380 0.000 703.920 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER ME3 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER ME2 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER ME1 ;
  RECT 639.620 0.000 643.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 626.600 0.000 630.140 1.120 ;
  LAYER ME3 ;
  RECT 626.600 0.000 630.140 1.120 ;
  LAYER ME2 ;
  RECT 626.600 0.000 630.140 1.120 ;
  LAYER ME1 ;
  RECT 626.600 0.000 630.140 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER ME3 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER ME2 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER ME1 ;
  RECT 604.900 0.000 608.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER ME3 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER ME2 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER ME1 ;
  RECT 596.220 0.000 599.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER ME3 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER ME2 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER ME1 ;
  RECT 587.540 0.000 591.080 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER ME3 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER ME2 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER ME1 ;
  RECT 578.860 0.000 582.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.680 0.000 465.220 1.120 ;
  LAYER ME3 ;
  RECT 461.680 0.000 465.220 1.120 ;
  LAYER ME2 ;
  RECT 461.680 0.000 465.220 1.120 ;
  LAYER ME1 ;
  RECT 461.680 0.000 465.220 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME3 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME2 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME1 ;
  RECT 453.000 0.000 456.540 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME3 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME2 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME1 ;
  RECT 444.320 0.000 447.860 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER ME3 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER ME2 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER ME1 ;
  RECT 435.640 0.000 439.180 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER ME3 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER ME2 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER ME1 ;
  RECT 422.620 0.000 426.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 400.920 0.000 404.460 1.120 ;
  LAYER ME3 ;
  RECT 400.920 0.000 404.460 1.120 ;
  LAYER ME2 ;
  RECT 400.920 0.000 404.460 1.120 ;
  LAYER ME1 ;
  RECT 400.920 0.000 404.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.160 0.000 343.700 1.120 ;
  LAYER ME3 ;
  RECT 340.160 0.000 343.700 1.120 ;
  LAYER ME2 ;
  RECT 340.160 0.000 343.700 1.120 ;
  LAYER ME1 ;
  RECT 340.160 0.000 343.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.480 0.000 335.020 1.120 ;
  LAYER ME3 ;
  RECT 331.480 0.000 335.020 1.120 ;
  LAYER ME2 ;
  RECT 331.480 0.000 335.020 1.120 ;
  LAYER ME1 ;
  RECT 331.480 0.000 335.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.800 0.000 326.340 1.120 ;
  LAYER ME3 ;
  RECT 322.800 0.000 326.340 1.120 ;
  LAYER ME2 ;
  RECT 322.800 0.000 326.340 1.120 ;
  LAYER ME1 ;
  RECT 322.800 0.000 326.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME3 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME2 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME1 ;
  RECT 309.780 0.000 313.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.460 0.000 291.000 1.120 ;
  LAYER ME3 ;
  RECT 287.460 0.000 291.000 1.120 ;
  LAYER ME2 ;
  RECT 287.460 0.000 291.000 1.120 ;
  LAYER ME1 ;
  RECT 287.460 0.000 291.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER ME3 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER ME2 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER ME1 ;
  RECT 278.780 0.000 282.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.680 0.000 217.220 1.120 ;
  LAYER ME3 ;
  RECT 213.680 0.000 217.220 1.120 ;
  LAYER ME2 ;
  RECT 213.680 0.000 217.220 1.120 ;
  LAYER ME1 ;
  RECT 213.680 0.000 217.220 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.000 0.000 208.540 1.120 ;
  LAYER ME3 ;
  RECT 205.000 0.000 208.540 1.120 ;
  LAYER ME2 ;
  RECT 205.000 0.000 208.540 1.120 ;
  LAYER ME1 ;
  RECT 205.000 0.000 208.540 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.300 0.000 186.840 1.120 ;
  LAYER ME3 ;
  RECT 183.300 0.000 186.840 1.120 ;
  LAYER ME2 ;
  RECT 183.300 0.000 186.840 1.120 ;
  LAYER ME1 ;
  RECT 183.300 0.000 186.840 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER ME3 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER ME2 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER ME1 ;
  RECT 170.280 0.000 173.820 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER ME3 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER ME2 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER ME1 ;
  RECT 161.600 0.000 165.140 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER ME3 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER ME2 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER ME1 ;
  RECT 152.920 0.000 156.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER ME3 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER ME2 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER ME1 ;
  RECT 57.440 0.000 60.980 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER ME3 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER ME2 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER ME1 ;
  RECT 48.760 0.000 52.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER ME3 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER ME2 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER ME1 ;
  RECT 40.080 0.000 43.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 1014.440 1376.260 1015.560 1379.500 ;
  LAYER ME3 ;
  RECT 1014.440 1376.260 1015.560 1379.500 ;
  LAYER ME2 ;
  RECT 1014.440 1376.260 1015.560 1379.500 ;
  LAYER ME1 ;
  RECT 1014.440 1376.260 1015.560 1379.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1368.420 1015.560 1371.660 ;
  LAYER ME3 ;
  RECT 1014.440 1368.420 1015.560 1371.660 ;
  LAYER ME2 ;
  RECT 1014.440 1368.420 1015.560 1371.660 ;
  LAYER ME1 ;
  RECT 1014.440 1368.420 1015.560 1371.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1360.580 1015.560 1363.820 ;
  LAYER ME3 ;
  RECT 1014.440 1360.580 1015.560 1363.820 ;
  LAYER ME2 ;
  RECT 1014.440 1360.580 1015.560 1363.820 ;
  LAYER ME1 ;
  RECT 1014.440 1360.580 1015.560 1363.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1352.740 1015.560 1355.980 ;
  LAYER ME3 ;
  RECT 1014.440 1352.740 1015.560 1355.980 ;
  LAYER ME2 ;
  RECT 1014.440 1352.740 1015.560 1355.980 ;
  LAYER ME1 ;
  RECT 1014.440 1352.740 1015.560 1355.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1344.900 1015.560 1348.140 ;
  LAYER ME3 ;
  RECT 1014.440 1344.900 1015.560 1348.140 ;
  LAYER ME2 ;
  RECT 1014.440 1344.900 1015.560 1348.140 ;
  LAYER ME1 ;
  RECT 1014.440 1344.900 1015.560 1348.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1305.700 1015.560 1308.940 ;
  LAYER ME3 ;
  RECT 1014.440 1305.700 1015.560 1308.940 ;
  LAYER ME2 ;
  RECT 1014.440 1305.700 1015.560 1308.940 ;
  LAYER ME1 ;
  RECT 1014.440 1305.700 1015.560 1308.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1297.860 1015.560 1301.100 ;
  LAYER ME3 ;
  RECT 1014.440 1297.860 1015.560 1301.100 ;
  LAYER ME2 ;
  RECT 1014.440 1297.860 1015.560 1301.100 ;
  LAYER ME1 ;
  RECT 1014.440 1297.860 1015.560 1301.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1290.020 1015.560 1293.260 ;
  LAYER ME3 ;
  RECT 1014.440 1290.020 1015.560 1293.260 ;
  LAYER ME2 ;
  RECT 1014.440 1290.020 1015.560 1293.260 ;
  LAYER ME1 ;
  RECT 1014.440 1290.020 1015.560 1293.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1282.180 1015.560 1285.420 ;
  LAYER ME3 ;
  RECT 1014.440 1282.180 1015.560 1285.420 ;
  LAYER ME2 ;
  RECT 1014.440 1282.180 1015.560 1285.420 ;
  LAYER ME1 ;
  RECT 1014.440 1282.180 1015.560 1285.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1274.340 1015.560 1277.580 ;
  LAYER ME3 ;
  RECT 1014.440 1274.340 1015.560 1277.580 ;
  LAYER ME2 ;
  RECT 1014.440 1274.340 1015.560 1277.580 ;
  LAYER ME1 ;
  RECT 1014.440 1274.340 1015.560 1277.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1266.500 1015.560 1269.740 ;
  LAYER ME3 ;
  RECT 1014.440 1266.500 1015.560 1269.740 ;
  LAYER ME2 ;
  RECT 1014.440 1266.500 1015.560 1269.740 ;
  LAYER ME1 ;
  RECT 1014.440 1266.500 1015.560 1269.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1227.300 1015.560 1230.540 ;
  LAYER ME3 ;
  RECT 1014.440 1227.300 1015.560 1230.540 ;
  LAYER ME2 ;
  RECT 1014.440 1227.300 1015.560 1230.540 ;
  LAYER ME1 ;
  RECT 1014.440 1227.300 1015.560 1230.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1219.460 1015.560 1222.700 ;
  LAYER ME3 ;
  RECT 1014.440 1219.460 1015.560 1222.700 ;
  LAYER ME2 ;
  RECT 1014.440 1219.460 1015.560 1222.700 ;
  LAYER ME1 ;
  RECT 1014.440 1219.460 1015.560 1222.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1211.620 1015.560 1214.860 ;
  LAYER ME3 ;
  RECT 1014.440 1211.620 1015.560 1214.860 ;
  LAYER ME2 ;
  RECT 1014.440 1211.620 1015.560 1214.860 ;
  LAYER ME1 ;
  RECT 1014.440 1211.620 1015.560 1214.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1203.780 1015.560 1207.020 ;
  LAYER ME3 ;
  RECT 1014.440 1203.780 1015.560 1207.020 ;
  LAYER ME2 ;
  RECT 1014.440 1203.780 1015.560 1207.020 ;
  LAYER ME1 ;
  RECT 1014.440 1203.780 1015.560 1207.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1195.940 1015.560 1199.180 ;
  LAYER ME3 ;
  RECT 1014.440 1195.940 1015.560 1199.180 ;
  LAYER ME2 ;
  RECT 1014.440 1195.940 1015.560 1199.180 ;
  LAYER ME1 ;
  RECT 1014.440 1195.940 1015.560 1199.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1188.100 1015.560 1191.340 ;
  LAYER ME3 ;
  RECT 1014.440 1188.100 1015.560 1191.340 ;
  LAYER ME2 ;
  RECT 1014.440 1188.100 1015.560 1191.340 ;
  LAYER ME1 ;
  RECT 1014.440 1188.100 1015.560 1191.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1148.900 1015.560 1152.140 ;
  LAYER ME3 ;
  RECT 1014.440 1148.900 1015.560 1152.140 ;
  LAYER ME2 ;
  RECT 1014.440 1148.900 1015.560 1152.140 ;
  LAYER ME1 ;
  RECT 1014.440 1148.900 1015.560 1152.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1141.060 1015.560 1144.300 ;
  LAYER ME3 ;
  RECT 1014.440 1141.060 1015.560 1144.300 ;
  LAYER ME2 ;
  RECT 1014.440 1141.060 1015.560 1144.300 ;
  LAYER ME1 ;
  RECT 1014.440 1141.060 1015.560 1144.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1133.220 1015.560 1136.460 ;
  LAYER ME3 ;
  RECT 1014.440 1133.220 1015.560 1136.460 ;
  LAYER ME2 ;
  RECT 1014.440 1133.220 1015.560 1136.460 ;
  LAYER ME1 ;
  RECT 1014.440 1133.220 1015.560 1136.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1125.380 1015.560 1128.620 ;
  LAYER ME3 ;
  RECT 1014.440 1125.380 1015.560 1128.620 ;
  LAYER ME2 ;
  RECT 1014.440 1125.380 1015.560 1128.620 ;
  LAYER ME1 ;
  RECT 1014.440 1125.380 1015.560 1128.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1117.540 1015.560 1120.780 ;
  LAYER ME3 ;
  RECT 1014.440 1117.540 1015.560 1120.780 ;
  LAYER ME2 ;
  RECT 1014.440 1117.540 1015.560 1120.780 ;
  LAYER ME1 ;
  RECT 1014.440 1117.540 1015.560 1120.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1109.700 1015.560 1112.940 ;
  LAYER ME3 ;
  RECT 1014.440 1109.700 1015.560 1112.940 ;
  LAYER ME2 ;
  RECT 1014.440 1109.700 1015.560 1112.940 ;
  LAYER ME1 ;
  RECT 1014.440 1109.700 1015.560 1112.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1070.500 1015.560 1073.740 ;
  LAYER ME3 ;
  RECT 1014.440 1070.500 1015.560 1073.740 ;
  LAYER ME2 ;
  RECT 1014.440 1070.500 1015.560 1073.740 ;
  LAYER ME1 ;
  RECT 1014.440 1070.500 1015.560 1073.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1062.660 1015.560 1065.900 ;
  LAYER ME3 ;
  RECT 1014.440 1062.660 1015.560 1065.900 ;
  LAYER ME2 ;
  RECT 1014.440 1062.660 1015.560 1065.900 ;
  LAYER ME1 ;
  RECT 1014.440 1062.660 1015.560 1065.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1054.820 1015.560 1058.060 ;
  LAYER ME3 ;
  RECT 1014.440 1054.820 1015.560 1058.060 ;
  LAYER ME2 ;
  RECT 1014.440 1054.820 1015.560 1058.060 ;
  LAYER ME1 ;
  RECT 1014.440 1054.820 1015.560 1058.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1046.980 1015.560 1050.220 ;
  LAYER ME3 ;
  RECT 1014.440 1046.980 1015.560 1050.220 ;
  LAYER ME2 ;
  RECT 1014.440 1046.980 1015.560 1050.220 ;
  LAYER ME1 ;
  RECT 1014.440 1046.980 1015.560 1050.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1039.140 1015.560 1042.380 ;
  LAYER ME3 ;
  RECT 1014.440 1039.140 1015.560 1042.380 ;
  LAYER ME2 ;
  RECT 1014.440 1039.140 1015.560 1042.380 ;
  LAYER ME1 ;
  RECT 1014.440 1039.140 1015.560 1042.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 1031.300 1015.560 1034.540 ;
  LAYER ME3 ;
  RECT 1014.440 1031.300 1015.560 1034.540 ;
  LAYER ME2 ;
  RECT 1014.440 1031.300 1015.560 1034.540 ;
  LAYER ME1 ;
  RECT 1014.440 1031.300 1015.560 1034.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 992.100 1015.560 995.340 ;
  LAYER ME3 ;
  RECT 1014.440 992.100 1015.560 995.340 ;
  LAYER ME2 ;
  RECT 1014.440 992.100 1015.560 995.340 ;
  LAYER ME1 ;
  RECT 1014.440 992.100 1015.560 995.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 984.260 1015.560 987.500 ;
  LAYER ME3 ;
  RECT 1014.440 984.260 1015.560 987.500 ;
  LAYER ME2 ;
  RECT 1014.440 984.260 1015.560 987.500 ;
  LAYER ME1 ;
  RECT 1014.440 984.260 1015.560 987.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 976.420 1015.560 979.660 ;
  LAYER ME3 ;
  RECT 1014.440 976.420 1015.560 979.660 ;
  LAYER ME2 ;
  RECT 1014.440 976.420 1015.560 979.660 ;
  LAYER ME1 ;
  RECT 1014.440 976.420 1015.560 979.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 968.580 1015.560 971.820 ;
  LAYER ME3 ;
  RECT 1014.440 968.580 1015.560 971.820 ;
  LAYER ME2 ;
  RECT 1014.440 968.580 1015.560 971.820 ;
  LAYER ME1 ;
  RECT 1014.440 968.580 1015.560 971.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 960.740 1015.560 963.980 ;
  LAYER ME3 ;
  RECT 1014.440 960.740 1015.560 963.980 ;
  LAYER ME2 ;
  RECT 1014.440 960.740 1015.560 963.980 ;
  LAYER ME1 ;
  RECT 1014.440 960.740 1015.560 963.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 952.900 1015.560 956.140 ;
  LAYER ME3 ;
  RECT 1014.440 952.900 1015.560 956.140 ;
  LAYER ME2 ;
  RECT 1014.440 952.900 1015.560 956.140 ;
  LAYER ME1 ;
  RECT 1014.440 952.900 1015.560 956.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 913.700 1015.560 916.940 ;
  LAYER ME3 ;
  RECT 1014.440 913.700 1015.560 916.940 ;
  LAYER ME2 ;
  RECT 1014.440 913.700 1015.560 916.940 ;
  LAYER ME1 ;
  RECT 1014.440 913.700 1015.560 916.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 905.860 1015.560 909.100 ;
  LAYER ME3 ;
  RECT 1014.440 905.860 1015.560 909.100 ;
  LAYER ME2 ;
  RECT 1014.440 905.860 1015.560 909.100 ;
  LAYER ME1 ;
  RECT 1014.440 905.860 1015.560 909.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 898.020 1015.560 901.260 ;
  LAYER ME3 ;
  RECT 1014.440 898.020 1015.560 901.260 ;
  LAYER ME2 ;
  RECT 1014.440 898.020 1015.560 901.260 ;
  LAYER ME1 ;
  RECT 1014.440 898.020 1015.560 901.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 890.180 1015.560 893.420 ;
  LAYER ME3 ;
  RECT 1014.440 890.180 1015.560 893.420 ;
  LAYER ME2 ;
  RECT 1014.440 890.180 1015.560 893.420 ;
  LAYER ME1 ;
  RECT 1014.440 890.180 1015.560 893.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 882.340 1015.560 885.580 ;
  LAYER ME3 ;
  RECT 1014.440 882.340 1015.560 885.580 ;
  LAYER ME2 ;
  RECT 1014.440 882.340 1015.560 885.580 ;
  LAYER ME1 ;
  RECT 1014.440 882.340 1015.560 885.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 874.500 1015.560 877.740 ;
  LAYER ME3 ;
  RECT 1014.440 874.500 1015.560 877.740 ;
  LAYER ME2 ;
  RECT 1014.440 874.500 1015.560 877.740 ;
  LAYER ME1 ;
  RECT 1014.440 874.500 1015.560 877.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 835.300 1015.560 838.540 ;
  LAYER ME3 ;
  RECT 1014.440 835.300 1015.560 838.540 ;
  LAYER ME2 ;
  RECT 1014.440 835.300 1015.560 838.540 ;
  LAYER ME1 ;
  RECT 1014.440 835.300 1015.560 838.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 827.460 1015.560 830.700 ;
  LAYER ME3 ;
  RECT 1014.440 827.460 1015.560 830.700 ;
  LAYER ME2 ;
  RECT 1014.440 827.460 1015.560 830.700 ;
  LAYER ME1 ;
  RECT 1014.440 827.460 1015.560 830.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 819.620 1015.560 822.860 ;
  LAYER ME3 ;
  RECT 1014.440 819.620 1015.560 822.860 ;
  LAYER ME2 ;
  RECT 1014.440 819.620 1015.560 822.860 ;
  LAYER ME1 ;
  RECT 1014.440 819.620 1015.560 822.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 811.780 1015.560 815.020 ;
  LAYER ME3 ;
  RECT 1014.440 811.780 1015.560 815.020 ;
  LAYER ME2 ;
  RECT 1014.440 811.780 1015.560 815.020 ;
  LAYER ME1 ;
  RECT 1014.440 811.780 1015.560 815.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 803.940 1015.560 807.180 ;
  LAYER ME3 ;
  RECT 1014.440 803.940 1015.560 807.180 ;
  LAYER ME2 ;
  RECT 1014.440 803.940 1015.560 807.180 ;
  LAYER ME1 ;
  RECT 1014.440 803.940 1015.560 807.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 796.100 1015.560 799.340 ;
  LAYER ME3 ;
  RECT 1014.440 796.100 1015.560 799.340 ;
  LAYER ME2 ;
  RECT 1014.440 796.100 1015.560 799.340 ;
  LAYER ME1 ;
  RECT 1014.440 796.100 1015.560 799.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 756.900 1015.560 760.140 ;
  LAYER ME3 ;
  RECT 1014.440 756.900 1015.560 760.140 ;
  LAYER ME2 ;
  RECT 1014.440 756.900 1015.560 760.140 ;
  LAYER ME1 ;
  RECT 1014.440 756.900 1015.560 760.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 749.060 1015.560 752.300 ;
  LAYER ME3 ;
  RECT 1014.440 749.060 1015.560 752.300 ;
  LAYER ME2 ;
  RECT 1014.440 749.060 1015.560 752.300 ;
  LAYER ME1 ;
  RECT 1014.440 749.060 1015.560 752.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 741.220 1015.560 744.460 ;
  LAYER ME3 ;
  RECT 1014.440 741.220 1015.560 744.460 ;
  LAYER ME2 ;
  RECT 1014.440 741.220 1015.560 744.460 ;
  LAYER ME1 ;
  RECT 1014.440 741.220 1015.560 744.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 733.380 1015.560 736.620 ;
  LAYER ME3 ;
  RECT 1014.440 733.380 1015.560 736.620 ;
  LAYER ME2 ;
  RECT 1014.440 733.380 1015.560 736.620 ;
  LAYER ME1 ;
  RECT 1014.440 733.380 1015.560 736.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 725.540 1015.560 728.780 ;
  LAYER ME3 ;
  RECT 1014.440 725.540 1015.560 728.780 ;
  LAYER ME2 ;
  RECT 1014.440 725.540 1015.560 728.780 ;
  LAYER ME1 ;
  RECT 1014.440 725.540 1015.560 728.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 717.700 1015.560 720.940 ;
  LAYER ME3 ;
  RECT 1014.440 717.700 1015.560 720.940 ;
  LAYER ME2 ;
  RECT 1014.440 717.700 1015.560 720.940 ;
  LAYER ME1 ;
  RECT 1014.440 717.700 1015.560 720.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 678.500 1015.560 681.740 ;
  LAYER ME3 ;
  RECT 1014.440 678.500 1015.560 681.740 ;
  LAYER ME2 ;
  RECT 1014.440 678.500 1015.560 681.740 ;
  LAYER ME1 ;
  RECT 1014.440 678.500 1015.560 681.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 670.660 1015.560 673.900 ;
  LAYER ME3 ;
  RECT 1014.440 670.660 1015.560 673.900 ;
  LAYER ME2 ;
  RECT 1014.440 670.660 1015.560 673.900 ;
  LAYER ME1 ;
  RECT 1014.440 670.660 1015.560 673.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 662.820 1015.560 666.060 ;
  LAYER ME3 ;
  RECT 1014.440 662.820 1015.560 666.060 ;
  LAYER ME2 ;
  RECT 1014.440 662.820 1015.560 666.060 ;
  LAYER ME1 ;
  RECT 1014.440 662.820 1015.560 666.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 654.980 1015.560 658.220 ;
  LAYER ME3 ;
  RECT 1014.440 654.980 1015.560 658.220 ;
  LAYER ME2 ;
  RECT 1014.440 654.980 1015.560 658.220 ;
  LAYER ME1 ;
  RECT 1014.440 654.980 1015.560 658.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 647.140 1015.560 650.380 ;
  LAYER ME3 ;
  RECT 1014.440 647.140 1015.560 650.380 ;
  LAYER ME2 ;
  RECT 1014.440 647.140 1015.560 650.380 ;
  LAYER ME1 ;
  RECT 1014.440 647.140 1015.560 650.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 639.300 1015.560 642.540 ;
  LAYER ME3 ;
  RECT 1014.440 639.300 1015.560 642.540 ;
  LAYER ME2 ;
  RECT 1014.440 639.300 1015.560 642.540 ;
  LAYER ME1 ;
  RECT 1014.440 639.300 1015.560 642.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 600.100 1015.560 603.340 ;
  LAYER ME3 ;
  RECT 1014.440 600.100 1015.560 603.340 ;
  LAYER ME2 ;
  RECT 1014.440 600.100 1015.560 603.340 ;
  LAYER ME1 ;
  RECT 1014.440 600.100 1015.560 603.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 592.260 1015.560 595.500 ;
  LAYER ME3 ;
  RECT 1014.440 592.260 1015.560 595.500 ;
  LAYER ME2 ;
  RECT 1014.440 592.260 1015.560 595.500 ;
  LAYER ME1 ;
  RECT 1014.440 592.260 1015.560 595.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 584.420 1015.560 587.660 ;
  LAYER ME3 ;
  RECT 1014.440 584.420 1015.560 587.660 ;
  LAYER ME2 ;
  RECT 1014.440 584.420 1015.560 587.660 ;
  LAYER ME1 ;
  RECT 1014.440 584.420 1015.560 587.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 576.580 1015.560 579.820 ;
  LAYER ME3 ;
  RECT 1014.440 576.580 1015.560 579.820 ;
  LAYER ME2 ;
  RECT 1014.440 576.580 1015.560 579.820 ;
  LAYER ME1 ;
  RECT 1014.440 576.580 1015.560 579.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 568.740 1015.560 571.980 ;
  LAYER ME3 ;
  RECT 1014.440 568.740 1015.560 571.980 ;
  LAYER ME2 ;
  RECT 1014.440 568.740 1015.560 571.980 ;
  LAYER ME1 ;
  RECT 1014.440 568.740 1015.560 571.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 560.900 1015.560 564.140 ;
  LAYER ME3 ;
  RECT 1014.440 560.900 1015.560 564.140 ;
  LAYER ME2 ;
  RECT 1014.440 560.900 1015.560 564.140 ;
  LAYER ME1 ;
  RECT 1014.440 560.900 1015.560 564.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 521.700 1015.560 524.940 ;
  LAYER ME3 ;
  RECT 1014.440 521.700 1015.560 524.940 ;
  LAYER ME2 ;
  RECT 1014.440 521.700 1015.560 524.940 ;
  LAYER ME1 ;
  RECT 1014.440 521.700 1015.560 524.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 513.860 1015.560 517.100 ;
  LAYER ME3 ;
  RECT 1014.440 513.860 1015.560 517.100 ;
  LAYER ME2 ;
  RECT 1014.440 513.860 1015.560 517.100 ;
  LAYER ME1 ;
  RECT 1014.440 513.860 1015.560 517.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 506.020 1015.560 509.260 ;
  LAYER ME3 ;
  RECT 1014.440 506.020 1015.560 509.260 ;
  LAYER ME2 ;
  RECT 1014.440 506.020 1015.560 509.260 ;
  LAYER ME1 ;
  RECT 1014.440 506.020 1015.560 509.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 498.180 1015.560 501.420 ;
  LAYER ME3 ;
  RECT 1014.440 498.180 1015.560 501.420 ;
  LAYER ME2 ;
  RECT 1014.440 498.180 1015.560 501.420 ;
  LAYER ME1 ;
  RECT 1014.440 498.180 1015.560 501.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 490.340 1015.560 493.580 ;
  LAYER ME3 ;
  RECT 1014.440 490.340 1015.560 493.580 ;
  LAYER ME2 ;
  RECT 1014.440 490.340 1015.560 493.580 ;
  LAYER ME1 ;
  RECT 1014.440 490.340 1015.560 493.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 482.500 1015.560 485.740 ;
  LAYER ME3 ;
  RECT 1014.440 482.500 1015.560 485.740 ;
  LAYER ME2 ;
  RECT 1014.440 482.500 1015.560 485.740 ;
  LAYER ME1 ;
  RECT 1014.440 482.500 1015.560 485.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 443.300 1015.560 446.540 ;
  LAYER ME3 ;
  RECT 1014.440 443.300 1015.560 446.540 ;
  LAYER ME2 ;
  RECT 1014.440 443.300 1015.560 446.540 ;
  LAYER ME1 ;
  RECT 1014.440 443.300 1015.560 446.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 435.460 1015.560 438.700 ;
  LAYER ME3 ;
  RECT 1014.440 435.460 1015.560 438.700 ;
  LAYER ME2 ;
  RECT 1014.440 435.460 1015.560 438.700 ;
  LAYER ME1 ;
  RECT 1014.440 435.460 1015.560 438.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 427.620 1015.560 430.860 ;
  LAYER ME3 ;
  RECT 1014.440 427.620 1015.560 430.860 ;
  LAYER ME2 ;
  RECT 1014.440 427.620 1015.560 430.860 ;
  LAYER ME1 ;
  RECT 1014.440 427.620 1015.560 430.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 419.780 1015.560 423.020 ;
  LAYER ME3 ;
  RECT 1014.440 419.780 1015.560 423.020 ;
  LAYER ME2 ;
  RECT 1014.440 419.780 1015.560 423.020 ;
  LAYER ME1 ;
  RECT 1014.440 419.780 1015.560 423.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 411.940 1015.560 415.180 ;
  LAYER ME3 ;
  RECT 1014.440 411.940 1015.560 415.180 ;
  LAYER ME2 ;
  RECT 1014.440 411.940 1015.560 415.180 ;
  LAYER ME1 ;
  RECT 1014.440 411.940 1015.560 415.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 404.100 1015.560 407.340 ;
  LAYER ME3 ;
  RECT 1014.440 404.100 1015.560 407.340 ;
  LAYER ME2 ;
  RECT 1014.440 404.100 1015.560 407.340 ;
  LAYER ME1 ;
  RECT 1014.440 404.100 1015.560 407.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 364.900 1015.560 368.140 ;
  LAYER ME3 ;
  RECT 1014.440 364.900 1015.560 368.140 ;
  LAYER ME2 ;
  RECT 1014.440 364.900 1015.560 368.140 ;
  LAYER ME1 ;
  RECT 1014.440 364.900 1015.560 368.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 357.060 1015.560 360.300 ;
  LAYER ME3 ;
  RECT 1014.440 357.060 1015.560 360.300 ;
  LAYER ME2 ;
  RECT 1014.440 357.060 1015.560 360.300 ;
  LAYER ME1 ;
  RECT 1014.440 357.060 1015.560 360.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 349.220 1015.560 352.460 ;
  LAYER ME3 ;
  RECT 1014.440 349.220 1015.560 352.460 ;
  LAYER ME2 ;
  RECT 1014.440 349.220 1015.560 352.460 ;
  LAYER ME1 ;
  RECT 1014.440 349.220 1015.560 352.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 341.380 1015.560 344.620 ;
  LAYER ME3 ;
  RECT 1014.440 341.380 1015.560 344.620 ;
  LAYER ME2 ;
  RECT 1014.440 341.380 1015.560 344.620 ;
  LAYER ME1 ;
  RECT 1014.440 341.380 1015.560 344.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 333.540 1015.560 336.780 ;
  LAYER ME3 ;
  RECT 1014.440 333.540 1015.560 336.780 ;
  LAYER ME2 ;
  RECT 1014.440 333.540 1015.560 336.780 ;
  LAYER ME1 ;
  RECT 1014.440 333.540 1015.560 336.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 325.700 1015.560 328.940 ;
  LAYER ME3 ;
  RECT 1014.440 325.700 1015.560 328.940 ;
  LAYER ME2 ;
  RECT 1014.440 325.700 1015.560 328.940 ;
  LAYER ME1 ;
  RECT 1014.440 325.700 1015.560 328.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 286.500 1015.560 289.740 ;
  LAYER ME3 ;
  RECT 1014.440 286.500 1015.560 289.740 ;
  LAYER ME2 ;
  RECT 1014.440 286.500 1015.560 289.740 ;
  LAYER ME1 ;
  RECT 1014.440 286.500 1015.560 289.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 278.660 1015.560 281.900 ;
  LAYER ME3 ;
  RECT 1014.440 278.660 1015.560 281.900 ;
  LAYER ME2 ;
  RECT 1014.440 278.660 1015.560 281.900 ;
  LAYER ME1 ;
  RECT 1014.440 278.660 1015.560 281.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 270.820 1015.560 274.060 ;
  LAYER ME3 ;
  RECT 1014.440 270.820 1015.560 274.060 ;
  LAYER ME2 ;
  RECT 1014.440 270.820 1015.560 274.060 ;
  LAYER ME1 ;
  RECT 1014.440 270.820 1015.560 274.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 262.980 1015.560 266.220 ;
  LAYER ME3 ;
  RECT 1014.440 262.980 1015.560 266.220 ;
  LAYER ME2 ;
  RECT 1014.440 262.980 1015.560 266.220 ;
  LAYER ME1 ;
  RECT 1014.440 262.980 1015.560 266.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 255.140 1015.560 258.380 ;
  LAYER ME3 ;
  RECT 1014.440 255.140 1015.560 258.380 ;
  LAYER ME2 ;
  RECT 1014.440 255.140 1015.560 258.380 ;
  LAYER ME1 ;
  RECT 1014.440 255.140 1015.560 258.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 247.300 1015.560 250.540 ;
  LAYER ME3 ;
  RECT 1014.440 247.300 1015.560 250.540 ;
  LAYER ME2 ;
  RECT 1014.440 247.300 1015.560 250.540 ;
  LAYER ME1 ;
  RECT 1014.440 247.300 1015.560 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 208.100 1015.560 211.340 ;
  LAYER ME3 ;
  RECT 1014.440 208.100 1015.560 211.340 ;
  LAYER ME2 ;
  RECT 1014.440 208.100 1015.560 211.340 ;
  LAYER ME1 ;
  RECT 1014.440 208.100 1015.560 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 200.260 1015.560 203.500 ;
  LAYER ME3 ;
  RECT 1014.440 200.260 1015.560 203.500 ;
  LAYER ME2 ;
  RECT 1014.440 200.260 1015.560 203.500 ;
  LAYER ME1 ;
  RECT 1014.440 200.260 1015.560 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 192.420 1015.560 195.660 ;
  LAYER ME3 ;
  RECT 1014.440 192.420 1015.560 195.660 ;
  LAYER ME2 ;
  RECT 1014.440 192.420 1015.560 195.660 ;
  LAYER ME1 ;
  RECT 1014.440 192.420 1015.560 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 184.580 1015.560 187.820 ;
  LAYER ME3 ;
  RECT 1014.440 184.580 1015.560 187.820 ;
  LAYER ME2 ;
  RECT 1014.440 184.580 1015.560 187.820 ;
  LAYER ME1 ;
  RECT 1014.440 184.580 1015.560 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 176.740 1015.560 179.980 ;
  LAYER ME3 ;
  RECT 1014.440 176.740 1015.560 179.980 ;
  LAYER ME2 ;
  RECT 1014.440 176.740 1015.560 179.980 ;
  LAYER ME1 ;
  RECT 1014.440 176.740 1015.560 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 168.900 1015.560 172.140 ;
  LAYER ME3 ;
  RECT 1014.440 168.900 1015.560 172.140 ;
  LAYER ME2 ;
  RECT 1014.440 168.900 1015.560 172.140 ;
  LAYER ME1 ;
  RECT 1014.440 168.900 1015.560 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 129.700 1015.560 132.940 ;
  LAYER ME3 ;
  RECT 1014.440 129.700 1015.560 132.940 ;
  LAYER ME2 ;
  RECT 1014.440 129.700 1015.560 132.940 ;
  LAYER ME1 ;
  RECT 1014.440 129.700 1015.560 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 121.860 1015.560 125.100 ;
  LAYER ME3 ;
  RECT 1014.440 121.860 1015.560 125.100 ;
  LAYER ME2 ;
  RECT 1014.440 121.860 1015.560 125.100 ;
  LAYER ME1 ;
  RECT 1014.440 121.860 1015.560 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 114.020 1015.560 117.260 ;
  LAYER ME3 ;
  RECT 1014.440 114.020 1015.560 117.260 ;
  LAYER ME2 ;
  RECT 1014.440 114.020 1015.560 117.260 ;
  LAYER ME1 ;
  RECT 1014.440 114.020 1015.560 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 106.180 1015.560 109.420 ;
  LAYER ME3 ;
  RECT 1014.440 106.180 1015.560 109.420 ;
  LAYER ME2 ;
  RECT 1014.440 106.180 1015.560 109.420 ;
  LAYER ME1 ;
  RECT 1014.440 106.180 1015.560 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 98.340 1015.560 101.580 ;
  LAYER ME3 ;
  RECT 1014.440 98.340 1015.560 101.580 ;
  LAYER ME2 ;
  RECT 1014.440 98.340 1015.560 101.580 ;
  LAYER ME1 ;
  RECT 1014.440 98.340 1015.560 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 90.500 1015.560 93.740 ;
  LAYER ME3 ;
  RECT 1014.440 90.500 1015.560 93.740 ;
  LAYER ME2 ;
  RECT 1014.440 90.500 1015.560 93.740 ;
  LAYER ME1 ;
  RECT 1014.440 90.500 1015.560 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 51.300 1015.560 54.540 ;
  LAYER ME3 ;
  RECT 1014.440 51.300 1015.560 54.540 ;
  LAYER ME2 ;
  RECT 1014.440 51.300 1015.560 54.540 ;
  LAYER ME1 ;
  RECT 1014.440 51.300 1015.560 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 43.460 1015.560 46.700 ;
  LAYER ME3 ;
  RECT 1014.440 43.460 1015.560 46.700 ;
  LAYER ME2 ;
  RECT 1014.440 43.460 1015.560 46.700 ;
  LAYER ME1 ;
  RECT 1014.440 43.460 1015.560 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 35.620 1015.560 38.860 ;
  LAYER ME3 ;
  RECT 1014.440 35.620 1015.560 38.860 ;
  LAYER ME2 ;
  RECT 1014.440 35.620 1015.560 38.860 ;
  LAYER ME1 ;
  RECT 1014.440 35.620 1015.560 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 27.780 1015.560 31.020 ;
  LAYER ME3 ;
  RECT 1014.440 27.780 1015.560 31.020 ;
  LAYER ME2 ;
  RECT 1014.440 27.780 1015.560 31.020 ;
  LAYER ME1 ;
  RECT 1014.440 27.780 1015.560 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 19.940 1015.560 23.180 ;
  LAYER ME3 ;
  RECT 1014.440 19.940 1015.560 23.180 ;
  LAYER ME2 ;
  RECT 1014.440 19.940 1015.560 23.180 ;
  LAYER ME1 ;
  RECT 1014.440 19.940 1015.560 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1014.440 12.100 1015.560 15.340 ;
  LAYER ME3 ;
  RECT 1014.440 12.100 1015.560 15.340 ;
  LAYER ME2 ;
  RECT 1014.440 12.100 1015.560 15.340 ;
  LAYER ME1 ;
  RECT 1014.440 12.100 1015.560 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1376.260 1.120 1379.500 ;
  LAYER ME3 ;
  RECT 0.000 1376.260 1.120 1379.500 ;
  LAYER ME2 ;
  RECT 0.000 1376.260 1.120 1379.500 ;
  LAYER ME1 ;
  RECT 0.000 1376.260 1.120 1379.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1368.420 1.120 1371.660 ;
  LAYER ME3 ;
  RECT 0.000 1368.420 1.120 1371.660 ;
  LAYER ME2 ;
  RECT 0.000 1368.420 1.120 1371.660 ;
  LAYER ME1 ;
  RECT 0.000 1368.420 1.120 1371.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1360.580 1.120 1363.820 ;
  LAYER ME3 ;
  RECT 0.000 1360.580 1.120 1363.820 ;
  LAYER ME2 ;
  RECT 0.000 1360.580 1.120 1363.820 ;
  LAYER ME1 ;
  RECT 0.000 1360.580 1.120 1363.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1352.740 1.120 1355.980 ;
  LAYER ME3 ;
  RECT 0.000 1352.740 1.120 1355.980 ;
  LAYER ME2 ;
  RECT 0.000 1352.740 1.120 1355.980 ;
  LAYER ME1 ;
  RECT 0.000 1352.740 1.120 1355.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1344.900 1.120 1348.140 ;
  LAYER ME3 ;
  RECT 0.000 1344.900 1.120 1348.140 ;
  LAYER ME2 ;
  RECT 0.000 1344.900 1.120 1348.140 ;
  LAYER ME1 ;
  RECT 0.000 1344.900 1.120 1348.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1305.700 1.120 1308.940 ;
  LAYER ME3 ;
  RECT 0.000 1305.700 1.120 1308.940 ;
  LAYER ME2 ;
  RECT 0.000 1305.700 1.120 1308.940 ;
  LAYER ME1 ;
  RECT 0.000 1305.700 1.120 1308.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1297.860 1.120 1301.100 ;
  LAYER ME3 ;
  RECT 0.000 1297.860 1.120 1301.100 ;
  LAYER ME2 ;
  RECT 0.000 1297.860 1.120 1301.100 ;
  LAYER ME1 ;
  RECT 0.000 1297.860 1.120 1301.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1290.020 1.120 1293.260 ;
  LAYER ME3 ;
  RECT 0.000 1290.020 1.120 1293.260 ;
  LAYER ME2 ;
  RECT 0.000 1290.020 1.120 1293.260 ;
  LAYER ME1 ;
  RECT 0.000 1290.020 1.120 1293.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1282.180 1.120 1285.420 ;
  LAYER ME3 ;
  RECT 0.000 1282.180 1.120 1285.420 ;
  LAYER ME2 ;
  RECT 0.000 1282.180 1.120 1285.420 ;
  LAYER ME1 ;
  RECT 0.000 1282.180 1.120 1285.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1274.340 1.120 1277.580 ;
  LAYER ME3 ;
  RECT 0.000 1274.340 1.120 1277.580 ;
  LAYER ME2 ;
  RECT 0.000 1274.340 1.120 1277.580 ;
  LAYER ME1 ;
  RECT 0.000 1274.340 1.120 1277.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1266.500 1.120 1269.740 ;
  LAYER ME3 ;
  RECT 0.000 1266.500 1.120 1269.740 ;
  LAYER ME2 ;
  RECT 0.000 1266.500 1.120 1269.740 ;
  LAYER ME1 ;
  RECT 0.000 1266.500 1.120 1269.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1227.300 1.120 1230.540 ;
  LAYER ME3 ;
  RECT 0.000 1227.300 1.120 1230.540 ;
  LAYER ME2 ;
  RECT 0.000 1227.300 1.120 1230.540 ;
  LAYER ME1 ;
  RECT 0.000 1227.300 1.120 1230.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1219.460 1.120 1222.700 ;
  LAYER ME3 ;
  RECT 0.000 1219.460 1.120 1222.700 ;
  LAYER ME2 ;
  RECT 0.000 1219.460 1.120 1222.700 ;
  LAYER ME1 ;
  RECT 0.000 1219.460 1.120 1222.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1211.620 1.120 1214.860 ;
  LAYER ME3 ;
  RECT 0.000 1211.620 1.120 1214.860 ;
  LAYER ME2 ;
  RECT 0.000 1211.620 1.120 1214.860 ;
  LAYER ME1 ;
  RECT 0.000 1211.620 1.120 1214.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1203.780 1.120 1207.020 ;
  LAYER ME3 ;
  RECT 0.000 1203.780 1.120 1207.020 ;
  LAYER ME2 ;
  RECT 0.000 1203.780 1.120 1207.020 ;
  LAYER ME1 ;
  RECT 0.000 1203.780 1.120 1207.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1195.940 1.120 1199.180 ;
  LAYER ME3 ;
  RECT 0.000 1195.940 1.120 1199.180 ;
  LAYER ME2 ;
  RECT 0.000 1195.940 1.120 1199.180 ;
  LAYER ME1 ;
  RECT 0.000 1195.940 1.120 1199.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1188.100 1.120 1191.340 ;
  LAYER ME3 ;
  RECT 0.000 1188.100 1.120 1191.340 ;
  LAYER ME2 ;
  RECT 0.000 1188.100 1.120 1191.340 ;
  LAYER ME1 ;
  RECT 0.000 1188.100 1.120 1191.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1148.900 1.120 1152.140 ;
  LAYER ME3 ;
  RECT 0.000 1148.900 1.120 1152.140 ;
  LAYER ME2 ;
  RECT 0.000 1148.900 1.120 1152.140 ;
  LAYER ME1 ;
  RECT 0.000 1148.900 1.120 1152.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1141.060 1.120 1144.300 ;
  LAYER ME3 ;
  RECT 0.000 1141.060 1.120 1144.300 ;
  LAYER ME2 ;
  RECT 0.000 1141.060 1.120 1144.300 ;
  LAYER ME1 ;
  RECT 0.000 1141.060 1.120 1144.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1133.220 1.120 1136.460 ;
  LAYER ME3 ;
  RECT 0.000 1133.220 1.120 1136.460 ;
  LAYER ME2 ;
  RECT 0.000 1133.220 1.120 1136.460 ;
  LAYER ME1 ;
  RECT 0.000 1133.220 1.120 1136.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1125.380 1.120 1128.620 ;
  LAYER ME3 ;
  RECT 0.000 1125.380 1.120 1128.620 ;
  LAYER ME2 ;
  RECT 0.000 1125.380 1.120 1128.620 ;
  LAYER ME1 ;
  RECT 0.000 1125.380 1.120 1128.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1117.540 1.120 1120.780 ;
  LAYER ME3 ;
  RECT 0.000 1117.540 1.120 1120.780 ;
  LAYER ME2 ;
  RECT 0.000 1117.540 1.120 1120.780 ;
  LAYER ME1 ;
  RECT 0.000 1117.540 1.120 1120.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1109.700 1.120 1112.940 ;
  LAYER ME3 ;
  RECT 0.000 1109.700 1.120 1112.940 ;
  LAYER ME2 ;
  RECT 0.000 1109.700 1.120 1112.940 ;
  LAYER ME1 ;
  RECT 0.000 1109.700 1.120 1112.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1070.500 1.120 1073.740 ;
  LAYER ME3 ;
  RECT 0.000 1070.500 1.120 1073.740 ;
  LAYER ME2 ;
  RECT 0.000 1070.500 1.120 1073.740 ;
  LAYER ME1 ;
  RECT 0.000 1070.500 1.120 1073.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER ME3 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER ME2 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER ME1 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER ME3 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER ME2 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER ME1 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER ME3 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER ME2 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER ME1 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER ME3 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER ME2 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER ME1 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER ME3 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER ME2 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER ME1 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER ME3 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER ME2 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER ME1 ;
  RECT 0.000 992.100 1.120 995.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER ME3 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER ME2 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER ME1 ;
  RECT 0.000 984.260 1.120 987.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER ME3 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER ME2 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER ME1 ;
  RECT 0.000 976.420 1.120 979.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER ME3 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER ME2 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER ME1 ;
  RECT 0.000 968.580 1.120 971.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER ME3 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER ME2 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER ME1 ;
  RECT 0.000 960.740 1.120 963.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER ME3 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER ME2 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER ME1 ;
  RECT 0.000 952.900 1.120 956.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER ME3 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER ME2 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER ME1 ;
  RECT 0.000 913.700 1.120 916.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER ME3 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER ME2 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER ME1 ;
  RECT 0.000 905.860 1.120 909.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER ME3 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER ME2 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER ME1 ;
  RECT 0.000 898.020 1.120 901.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER ME3 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER ME2 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER ME1 ;
  RECT 0.000 890.180 1.120 893.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER ME3 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER ME2 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER ME1 ;
  RECT 0.000 882.340 1.120 885.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER ME3 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER ME2 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER ME1 ;
  RECT 0.000 874.500 1.120 877.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER ME3 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER ME2 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER ME1 ;
  RECT 0.000 835.300 1.120 838.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER ME3 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER ME2 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER ME1 ;
  RECT 0.000 827.460 1.120 830.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER ME3 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER ME2 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER ME1 ;
  RECT 0.000 819.620 1.120 822.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER ME3 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER ME2 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER ME1 ;
  RECT 0.000 811.780 1.120 815.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER ME3 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER ME2 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER ME1 ;
  RECT 0.000 803.940 1.120 807.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER ME3 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER ME2 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER ME1 ;
  RECT 0.000 796.100 1.120 799.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER ME3 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER ME2 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER ME1 ;
  RECT 0.000 756.900 1.120 760.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER ME3 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER ME2 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER ME1 ;
  RECT 0.000 749.060 1.120 752.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER ME3 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER ME2 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER ME1 ;
  RECT 0.000 741.220 1.120 744.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER ME3 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER ME2 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER ME1 ;
  RECT 0.000 733.380 1.120 736.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER ME3 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER ME2 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER ME1 ;
  RECT 0.000 725.540 1.120 728.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER ME3 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER ME2 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER ME1 ;
  RECT 0.000 717.700 1.120 720.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER ME3 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER ME2 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER ME1 ;
  RECT 0.000 678.500 1.120 681.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER ME3 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER ME2 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER ME1 ;
  RECT 0.000 670.660 1.120 673.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER ME3 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER ME2 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER ME1 ;
  RECT 0.000 662.820 1.120 666.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER ME3 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER ME2 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER ME1 ;
  RECT 0.000 654.980 1.120 658.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER ME3 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER ME2 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER ME1 ;
  RECT 0.000 647.140 1.120 650.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER ME3 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER ME2 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER ME1 ;
  RECT 0.000 639.300 1.120 642.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER ME3 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER ME2 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER ME1 ;
  RECT 0.000 600.100 1.120 603.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER ME3 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER ME2 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER ME1 ;
  RECT 0.000 592.260 1.120 595.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER ME3 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER ME2 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER ME1 ;
  RECT 0.000 584.420 1.120 587.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER ME3 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER ME2 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER ME1 ;
  RECT 0.000 576.580 1.120 579.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER ME3 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER ME2 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER ME1 ;
  RECT 0.000 568.740 1.120 571.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER ME3 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER ME2 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER ME1 ;
  RECT 0.000 560.900 1.120 564.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER ME3 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER ME2 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER ME1 ;
  RECT 0.000 521.700 1.120 524.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER ME3 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER ME2 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER ME1 ;
  RECT 0.000 513.860 1.120 517.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER ME3 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER ME2 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER ME1 ;
  RECT 0.000 506.020 1.120 509.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER ME3 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER ME2 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER ME1 ;
  RECT 0.000 498.180 1.120 501.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER ME3 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER ME2 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER ME1 ;
  RECT 0.000 490.340 1.120 493.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER ME3 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER ME2 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER ME1 ;
  RECT 0.000 482.500 1.120 485.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER ME3 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER ME2 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER ME1 ;
  RECT 0.000 443.300 1.120 446.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER ME3 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER ME2 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER ME1 ;
  RECT 0.000 435.460 1.120 438.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER ME3 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER ME2 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER ME1 ;
  RECT 0.000 427.620 1.120 430.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER ME3 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER ME2 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER ME1 ;
  RECT 0.000 419.780 1.120 423.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER ME3 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER ME2 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER ME1 ;
  RECT 0.000 411.940 1.120 415.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER ME3 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER ME2 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER ME1 ;
  RECT 0.000 404.100 1.120 407.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER ME3 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER ME2 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER ME1 ;
  RECT 0.000 364.900 1.120 368.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER ME3 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER ME2 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER ME1 ;
  RECT 0.000 357.060 1.120 360.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER ME3 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER ME2 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER ME1 ;
  RECT 0.000 349.220 1.120 352.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER ME3 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER ME2 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER ME1 ;
  RECT 0.000 341.380 1.120 344.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER ME3 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER ME2 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER ME1 ;
  RECT 0.000 333.540 1.120 336.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER ME3 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER ME2 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER ME1 ;
  RECT 0.000 325.700 1.120 328.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER ME3 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER ME2 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER ME1 ;
  RECT 0.000 286.500 1.120 289.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1001.700 1390.480 1005.240 1391.600 ;
  LAYER ME3 ;
  RECT 1001.700 1390.480 1005.240 1391.600 ;
  LAYER ME2 ;
  RECT 1001.700 1390.480 1005.240 1391.600 ;
  LAYER ME1 ;
  RECT 1001.700 1390.480 1005.240 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.020 1390.480 996.560 1391.600 ;
  LAYER ME3 ;
  RECT 993.020 1390.480 996.560 1391.600 ;
  LAYER ME2 ;
  RECT 993.020 1390.480 996.560 1391.600 ;
  LAYER ME1 ;
  RECT 993.020 1390.480 996.560 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 984.340 1390.480 987.880 1391.600 ;
  LAYER ME3 ;
  RECT 984.340 1390.480 987.880 1391.600 ;
  LAYER ME2 ;
  RECT 984.340 1390.480 987.880 1391.600 ;
  LAYER ME1 ;
  RECT 984.340 1390.480 987.880 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 975.660 1390.480 979.200 1391.600 ;
  LAYER ME3 ;
  RECT 975.660 1390.480 979.200 1391.600 ;
  LAYER ME2 ;
  RECT 975.660 1390.480 979.200 1391.600 ;
  LAYER ME1 ;
  RECT 975.660 1390.480 979.200 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 966.980 1390.480 970.520 1391.600 ;
  LAYER ME3 ;
  RECT 966.980 1390.480 970.520 1391.600 ;
  LAYER ME2 ;
  RECT 966.980 1390.480 970.520 1391.600 ;
  LAYER ME1 ;
  RECT 966.980 1390.480 970.520 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 923.580 1390.480 927.120 1391.600 ;
  LAYER ME3 ;
  RECT 923.580 1390.480 927.120 1391.600 ;
  LAYER ME2 ;
  RECT 923.580 1390.480 927.120 1391.600 ;
  LAYER ME1 ;
  RECT 923.580 1390.480 927.120 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 914.900 1390.480 918.440 1391.600 ;
  LAYER ME3 ;
  RECT 914.900 1390.480 918.440 1391.600 ;
  LAYER ME2 ;
  RECT 914.900 1390.480 918.440 1391.600 ;
  LAYER ME1 ;
  RECT 914.900 1390.480 918.440 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 906.220 1390.480 909.760 1391.600 ;
  LAYER ME3 ;
  RECT 906.220 1390.480 909.760 1391.600 ;
  LAYER ME2 ;
  RECT 906.220 1390.480 909.760 1391.600 ;
  LAYER ME1 ;
  RECT 906.220 1390.480 909.760 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 897.540 1390.480 901.080 1391.600 ;
  LAYER ME3 ;
  RECT 897.540 1390.480 901.080 1391.600 ;
  LAYER ME2 ;
  RECT 897.540 1390.480 901.080 1391.600 ;
  LAYER ME1 ;
  RECT 897.540 1390.480 901.080 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 888.860 1390.480 892.400 1391.600 ;
  LAYER ME3 ;
  RECT 888.860 1390.480 892.400 1391.600 ;
  LAYER ME2 ;
  RECT 888.860 1390.480 892.400 1391.600 ;
  LAYER ME1 ;
  RECT 888.860 1390.480 892.400 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 880.180 1390.480 883.720 1391.600 ;
  LAYER ME3 ;
  RECT 880.180 1390.480 883.720 1391.600 ;
  LAYER ME2 ;
  RECT 880.180 1390.480 883.720 1391.600 ;
  LAYER ME1 ;
  RECT 880.180 1390.480 883.720 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 836.780 1390.480 840.320 1391.600 ;
  LAYER ME3 ;
  RECT 836.780 1390.480 840.320 1391.600 ;
  LAYER ME2 ;
  RECT 836.780 1390.480 840.320 1391.600 ;
  LAYER ME1 ;
  RECT 836.780 1390.480 840.320 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 828.100 1390.480 831.640 1391.600 ;
  LAYER ME3 ;
  RECT 828.100 1390.480 831.640 1391.600 ;
  LAYER ME2 ;
  RECT 828.100 1390.480 831.640 1391.600 ;
  LAYER ME1 ;
  RECT 828.100 1390.480 831.640 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 819.420 1390.480 822.960 1391.600 ;
  LAYER ME3 ;
  RECT 819.420 1390.480 822.960 1391.600 ;
  LAYER ME2 ;
  RECT 819.420 1390.480 822.960 1391.600 ;
  LAYER ME1 ;
  RECT 819.420 1390.480 822.960 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 810.740 1390.480 814.280 1391.600 ;
  LAYER ME3 ;
  RECT 810.740 1390.480 814.280 1391.600 ;
  LAYER ME2 ;
  RECT 810.740 1390.480 814.280 1391.600 ;
  LAYER ME1 ;
  RECT 810.740 1390.480 814.280 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 802.060 1390.480 805.600 1391.600 ;
  LAYER ME3 ;
  RECT 802.060 1390.480 805.600 1391.600 ;
  LAYER ME2 ;
  RECT 802.060 1390.480 805.600 1391.600 ;
  LAYER ME1 ;
  RECT 802.060 1390.480 805.600 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 793.380 1390.480 796.920 1391.600 ;
  LAYER ME3 ;
  RECT 793.380 1390.480 796.920 1391.600 ;
  LAYER ME2 ;
  RECT 793.380 1390.480 796.920 1391.600 ;
  LAYER ME1 ;
  RECT 793.380 1390.480 796.920 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 749.980 1390.480 753.520 1391.600 ;
  LAYER ME3 ;
  RECT 749.980 1390.480 753.520 1391.600 ;
  LAYER ME2 ;
  RECT 749.980 1390.480 753.520 1391.600 ;
  LAYER ME1 ;
  RECT 749.980 1390.480 753.520 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 741.300 1390.480 744.840 1391.600 ;
  LAYER ME3 ;
  RECT 741.300 1390.480 744.840 1391.600 ;
  LAYER ME2 ;
  RECT 741.300 1390.480 744.840 1391.600 ;
  LAYER ME1 ;
  RECT 741.300 1390.480 744.840 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 732.620 1390.480 736.160 1391.600 ;
  LAYER ME3 ;
  RECT 732.620 1390.480 736.160 1391.600 ;
  LAYER ME2 ;
  RECT 732.620 1390.480 736.160 1391.600 ;
  LAYER ME1 ;
  RECT 732.620 1390.480 736.160 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 723.940 1390.480 727.480 1391.600 ;
  LAYER ME3 ;
  RECT 723.940 1390.480 727.480 1391.600 ;
  LAYER ME2 ;
  RECT 723.940 1390.480 727.480 1391.600 ;
  LAYER ME1 ;
  RECT 723.940 1390.480 727.480 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 715.260 1390.480 718.800 1391.600 ;
  LAYER ME3 ;
  RECT 715.260 1390.480 718.800 1391.600 ;
  LAYER ME2 ;
  RECT 715.260 1390.480 718.800 1391.600 ;
  LAYER ME1 ;
  RECT 715.260 1390.480 718.800 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 706.580 1390.480 710.120 1391.600 ;
  LAYER ME3 ;
  RECT 706.580 1390.480 710.120 1391.600 ;
  LAYER ME2 ;
  RECT 706.580 1390.480 710.120 1391.600 ;
  LAYER ME1 ;
  RECT 706.580 1390.480 710.120 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 663.180 1390.480 666.720 1391.600 ;
  LAYER ME3 ;
  RECT 663.180 1390.480 666.720 1391.600 ;
  LAYER ME2 ;
  RECT 663.180 1390.480 666.720 1391.600 ;
  LAYER ME1 ;
  RECT 663.180 1390.480 666.720 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.500 1390.480 658.040 1391.600 ;
  LAYER ME3 ;
  RECT 654.500 1390.480 658.040 1391.600 ;
  LAYER ME2 ;
  RECT 654.500 1390.480 658.040 1391.600 ;
  LAYER ME1 ;
  RECT 654.500 1390.480 658.040 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 645.820 1390.480 649.360 1391.600 ;
  LAYER ME3 ;
  RECT 645.820 1390.480 649.360 1391.600 ;
  LAYER ME2 ;
  RECT 645.820 1390.480 649.360 1391.600 ;
  LAYER ME1 ;
  RECT 645.820 1390.480 649.360 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 637.140 1390.480 640.680 1391.600 ;
  LAYER ME3 ;
  RECT 637.140 1390.480 640.680 1391.600 ;
  LAYER ME2 ;
  RECT 637.140 1390.480 640.680 1391.600 ;
  LAYER ME1 ;
  RECT 637.140 1390.480 640.680 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 628.460 1390.480 632.000 1391.600 ;
  LAYER ME3 ;
  RECT 628.460 1390.480 632.000 1391.600 ;
  LAYER ME2 ;
  RECT 628.460 1390.480 632.000 1391.600 ;
  LAYER ME1 ;
  RECT 628.460 1390.480 632.000 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 619.780 1390.480 623.320 1391.600 ;
  LAYER ME3 ;
  RECT 619.780 1390.480 623.320 1391.600 ;
  LAYER ME2 ;
  RECT 619.780 1390.480 623.320 1391.600 ;
  LAYER ME1 ;
  RECT 619.780 1390.480 623.320 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 576.380 1390.480 579.920 1391.600 ;
  LAYER ME3 ;
  RECT 576.380 1390.480 579.920 1391.600 ;
  LAYER ME2 ;
  RECT 576.380 1390.480 579.920 1391.600 ;
  LAYER ME1 ;
  RECT 576.380 1390.480 579.920 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 567.700 1390.480 571.240 1391.600 ;
  LAYER ME3 ;
  RECT 567.700 1390.480 571.240 1391.600 ;
  LAYER ME2 ;
  RECT 567.700 1390.480 571.240 1391.600 ;
  LAYER ME1 ;
  RECT 567.700 1390.480 571.240 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 559.020 1390.480 562.560 1391.600 ;
  LAYER ME3 ;
  RECT 559.020 1390.480 562.560 1391.600 ;
  LAYER ME2 ;
  RECT 559.020 1390.480 562.560 1391.600 ;
  LAYER ME1 ;
  RECT 559.020 1390.480 562.560 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.340 1390.480 553.880 1391.600 ;
  LAYER ME3 ;
  RECT 550.340 1390.480 553.880 1391.600 ;
  LAYER ME2 ;
  RECT 550.340 1390.480 553.880 1391.600 ;
  LAYER ME1 ;
  RECT 550.340 1390.480 553.880 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.660 1390.480 545.200 1391.600 ;
  LAYER ME3 ;
  RECT 541.660 1390.480 545.200 1391.600 ;
  LAYER ME2 ;
  RECT 541.660 1390.480 545.200 1391.600 ;
  LAYER ME1 ;
  RECT 541.660 1390.480 545.200 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.980 1390.480 536.520 1391.600 ;
  LAYER ME3 ;
  RECT 532.980 1390.480 536.520 1391.600 ;
  LAYER ME2 ;
  RECT 532.980 1390.480 536.520 1391.600 ;
  LAYER ME1 ;
  RECT 532.980 1390.480 536.520 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.580 1390.480 493.120 1391.600 ;
  LAYER ME3 ;
  RECT 489.580 1390.480 493.120 1391.600 ;
  LAYER ME2 ;
  RECT 489.580 1390.480 493.120 1391.600 ;
  LAYER ME1 ;
  RECT 489.580 1390.480 493.120 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.900 1390.480 484.440 1391.600 ;
  LAYER ME3 ;
  RECT 480.900 1390.480 484.440 1391.600 ;
  LAYER ME2 ;
  RECT 480.900 1390.480 484.440 1391.600 ;
  LAYER ME1 ;
  RECT 480.900 1390.480 484.440 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 1390.480 475.760 1391.600 ;
  LAYER ME3 ;
  RECT 472.220 1390.480 475.760 1391.600 ;
  LAYER ME2 ;
  RECT 472.220 1390.480 475.760 1391.600 ;
  LAYER ME1 ;
  RECT 472.220 1390.480 475.760 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.540 1390.480 467.080 1391.600 ;
  LAYER ME3 ;
  RECT 463.540 1390.480 467.080 1391.600 ;
  LAYER ME2 ;
  RECT 463.540 1390.480 467.080 1391.600 ;
  LAYER ME1 ;
  RECT 463.540 1390.480 467.080 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.860 1390.480 458.400 1391.600 ;
  LAYER ME3 ;
  RECT 454.860 1390.480 458.400 1391.600 ;
  LAYER ME2 ;
  RECT 454.860 1390.480 458.400 1391.600 ;
  LAYER ME1 ;
  RECT 454.860 1390.480 458.400 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.180 1390.480 449.720 1391.600 ;
  LAYER ME3 ;
  RECT 446.180 1390.480 449.720 1391.600 ;
  LAYER ME2 ;
  RECT 446.180 1390.480 449.720 1391.600 ;
  LAYER ME1 ;
  RECT 446.180 1390.480 449.720 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 1390.480 406.320 1391.600 ;
  LAYER ME3 ;
  RECT 402.780 1390.480 406.320 1391.600 ;
  LAYER ME2 ;
  RECT 402.780 1390.480 406.320 1391.600 ;
  LAYER ME1 ;
  RECT 402.780 1390.480 406.320 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.100 1390.480 397.640 1391.600 ;
  LAYER ME3 ;
  RECT 394.100 1390.480 397.640 1391.600 ;
  LAYER ME2 ;
  RECT 394.100 1390.480 397.640 1391.600 ;
  LAYER ME1 ;
  RECT 394.100 1390.480 397.640 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.420 1390.480 388.960 1391.600 ;
  LAYER ME3 ;
  RECT 385.420 1390.480 388.960 1391.600 ;
  LAYER ME2 ;
  RECT 385.420 1390.480 388.960 1391.600 ;
  LAYER ME1 ;
  RECT 385.420 1390.480 388.960 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.740 1390.480 380.280 1391.600 ;
  LAYER ME3 ;
  RECT 376.740 1390.480 380.280 1391.600 ;
  LAYER ME2 ;
  RECT 376.740 1390.480 380.280 1391.600 ;
  LAYER ME1 ;
  RECT 376.740 1390.480 380.280 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.060 1390.480 371.600 1391.600 ;
  LAYER ME3 ;
  RECT 368.060 1390.480 371.600 1391.600 ;
  LAYER ME2 ;
  RECT 368.060 1390.480 371.600 1391.600 ;
  LAYER ME1 ;
  RECT 368.060 1390.480 371.600 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.380 1390.480 362.920 1391.600 ;
  LAYER ME3 ;
  RECT 359.380 1390.480 362.920 1391.600 ;
  LAYER ME2 ;
  RECT 359.380 1390.480 362.920 1391.600 ;
  LAYER ME1 ;
  RECT 359.380 1390.480 362.920 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.980 1390.480 319.520 1391.600 ;
  LAYER ME3 ;
  RECT 315.980 1390.480 319.520 1391.600 ;
  LAYER ME2 ;
  RECT 315.980 1390.480 319.520 1391.600 ;
  LAYER ME1 ;
  RECT 315.980 1390.480 319.520 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 1390.480 310.840 1391.600 ;
  LAYER ME3 ;
  RECT 307.300 1390.480 310.840 1391.600 ;
  LAYER ME2 ;
  RECT 307.300 1390.480 310.840 1391.600 ;
  LAYER ME1 ;
  RECT 307.300 1390.480 310.840 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 1390.480 302.160 1391.600 ;
  LAYER ME3 ;
  RECT 298.620 1390.480 302.160 1391.600 ;
  LAYER ME2 ;
  RECT 298.620 1390.480 302.160 1391.600 ;
  LAYER ME1 ;
  RECT 298.620 1390.480 302.160 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 1390.480 293.480 1391.600 ;
  LAYER ME3 ;
  RECT 289.940 1390.480 293.480 1391.600 ;
  LAYER ME2 ;
  RECT 289.940 1390.480 293.480 1391.600 ;
  LAYER ME1 ;
  RECT 289.940 1390.480 293.480 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 1390.480 284.800 1391.600 ;
  LAYER ME3 ;
  RECT 281.260 1390.480 284.800 1391.600 ;
  LAYER ME2 ;
  RECT 281.260 1390.480 284.800 1391.600 ;
  LAYER ME1 ;
  RECT 281.260 1390.480 284.800 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 1390.480 276.120 1391.600 ;
  LAYER ME3 ;
  RECT 272.580 1390.480 276.120 1391.600 ;
  LAYER ME2 ;
  RECT 272.580 1390.480 276.120 1391.600 ;
  LAYER ME1 ;
  RECT 272.580 1390.480 276.120 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 1390.480 232.720 1391.600 ;
  LAYER ME3 ;
  RECT 229.180 1390.480 232.720 1391.600 ;
  LAYER ME2 ;
  RECT 229.180 1390.480 232.720 1391.600 ;
  LAYER ME1 ;
  RECT 229.180 1390.480 232.720 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 1390.480 224.040 1391.600 ;
  LAYER ME3 ;
  RECT 220.500 1390.480 224.040 1391.600 ;
  LAYER ME2 ;
  RECT 220.500 1390.480 224.040 1391.600 ;
  LAYER ME1 ;
  RECT 220.500 1390.480 224.040 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 1390.480 215.360 1391.600 ;
  LAYER ME3 ;
  RECT 211.820 1390.480 215.360 1391.600 ;
  LAYER ME2 ;
  RECT 211.820 1390.480 215.360 1391.600 ;
  LAYER ME1 ;
  RECT 211.820 1390.480 215.360 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 1390.480 206.680 1391.600 ;
  LAYER ME3 ;
  RECT 203.140 1390.480 206.680 1391.600 ;
  LAYER ME2 ;
  RECT 203.140 1390.480 206.680 1391.600 ;
  LAYER ME1 ;
  RECT 203.140 1390.480 206.680 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 1390.480 198.000 1391.600 ;
  LAYER ME3 ;
  RECT 194.460 1390.480 198.000 1391.600 ;
  LAYER ME2 ;
  RECT 194.460 1390.480 198.000 1391.600 ;
  LAYER ME1 ;
  RECT 194.460 1390.480 198.000 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 1390.480 189.320 1391.600 ;
  LAYER ME3 ;
  RECT 185.780 1390.480 189.320 1391.600 ;
  LAYER ME2 ;
  RECT 185.780 1390.480 189.320 1391.600 ;
  LAYER ME1 ;
  RECT 185.780 1390.480 189.320 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 1390.480 145.920 1391.600 ;
  LAYER ME3 ;
  RECT 142.380 1390.480 145.920 1391.600 ;
  LAYER ME2 ;
  RECT 142.380 1390.480 145.920 1391.600 ;
  LAYER ME1 ;
  RECT 142.380 1390.480 145.920 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 1390.480 137.240 1391.600 ;
  LAYER ME3 ;
  RECT 133.700 1390.480 137.240 1391.600 ;
  LAYER ME2 ;
  RECT 133.700 1390.480 137.240 1391.600 ;
  LAYER ME1 ;
  RECT 133.700 1390.480 137.240 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 1390.480 128.560 1391.600 ;
  LAYER ME3 ;
  RECT 125.020 1390.480 128.560 1391.600 ;
  LAYER ME2 ;
  RECT 125.020 1390.480 128.560 1391.600 ;
  LAYER ME1 ;
  RECT 125.020 1390.480 128.560 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 1390.480 119.880 1391.600 ;
  LAYER ME3 ;
  RECT 116.340 1390.480 119.880 1391.600 ;
  LAYER ME2 ;
  RECT 116.340 1390.480 119.880 1391.600 ;
  LAYER ME1 ;
  RECT 116.340 1390.480 119.880 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 1390.480 111.200 1391.600 ;
  LAYER ME3 ;
  RECT 107.660 1390.480 111.200 1391.600 ;
  LAYER ME2 ;
  RECT 107.660 1390.480 111.200 1391.600 ;
  LAYER ME1 ;
  RECT 107.660 1390.480 111.200 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 1390.480 102.520 1391.600 ;
  LAYER ME3 ;
  RECT 98.980 1390.480 102.520 1391.600 ;
  LAYER ME2 ;
  RECT 98.980 1390.480 102.520 1391.600 ;
  LAYER ME1 ;
  RECT 98.980 1390.480 102.520 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 1390.480 59.120 1391.600 ;
  LAYER ME3 ;
  RECT 55.580 1390.480 59.120 1391.600 ;
  LAYER ME2 ;
  RECT 55.580 1390.480 59.120 1391.600 ;
  LAYER ME1 ;
  RECT 55.580 1390.480 59.120 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 1390.480 50.440 1391.600 ;
  LAYER ME3 ;
  RECT 46.900 1390.480 50.440 1391.600 ;
  LAYER ME2 ;
  RECT 46.900 1390.480 50.440 1391.600 ;
  LAYER ME1 ;
  RECT 46.900 1390.480 50.440 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 1390.480 41.760 1391.600 ;
  LAYER ME3 ;
  RECT 38.220 1390.480 41.760 1391.600 ;
  LAYER ME2 ;
  RECT 38.220 1390.480 41.760 1391.600 ;
  LAYER ME1 ;
  RECT 38.220 1390.480 41.760 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 1390.480 33.080 1391.600 ;
  LAYER ME3 ;
  RECT 29.540 1390.480 33.080 1391.600 ;
  LAYER ME2 ;
  RECT 29.540 1390.480 33.080 1391.600 ;
  LAYER ME1 ;
  RECT 29.540 1390.480 33.080 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 1390.480 24.400 1391.600 ;
  LAYER ME3 ;
  RECT 20.860 1390.480 24.400 1391.600 ;
  LAYER ME2 ;
  RECT 20.860 1390.480 24.400 1391.600 ;
  LAYER ME1 ;
  RECT 20.860 1390.480 24.400 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 1390.480 15.720 1391.600 ;
  LAYER ME3 ;
  RECT 12.180 1390.480 15.720 1391.600 ;
  LAYER ME2 ;
  RECT 12.180 1390.480 15.720 1391.600 ;
  LAYER ME1 ;
  RECT 12.180 1390.480 15.720 1391.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER ME3 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER ME2 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER ME1 ;
  RECT 996.120 0.000 999.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 987.440 0.000 990.980 1.120 ;
  LAYER ME3 ;
  RECT 987.440 0.000 990.980 1.120 ;
  LAYER ME2 ;
  RECT 987.440 0.000 990.980 1.120 ;
  LAYER ME1 ;
  RECT 987.440 0.000 990.980 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 978.760 0.000 982.300 1.120 ;
  LAYER ME3 ;
  RECT 978.760 0.000 982.300 1.120 ;
  LAYER ME2 ;
  RECT 978.760 0.000 982.300 1.120 ;
  LAYER ME1 ;
  RECT 978.760 0.000 982.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 965.740 0.000 969.280 1.120 ;
  LAYER ME3 ;
  RECT 965.740 0.000 969.280 1.120 ;
  LAYER ME2 ;
  RECT 965.740 0.000 969.280 1.120 ;
  LAYER ME1 ;
  RECT 965.740 0.000 969.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 896.300 0.000 899.840 1.120 ;
  LAYER ME3 ;
  RECT 896.300 0.000 899.840 1.120 ;
  LAYER ME2 ;
  RECT 896.300 0.000 899.840 1.120 ;
  LAYER ME1 ;
  RECT 896.300 0.000 899.840 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER ME3 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER ME2 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER ME1 ;
  RECT 883.280 0.000 886.820 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER ME3 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER ME2 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER ME1 ;
  RECT 874.600 0.000 878.140 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER ME3 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER ME2 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER ME1 ;
  RECT 865.920 0.000 869.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER ME3 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER ME2 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER ME1 ;
  RECT 852.900 0.000 856.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER ME3 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER ME2 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER ME1 ;
  RECT 830.580 0.000 834.120 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER ME3 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER ME2 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER ME1 ;
  RECT 765.480 0.000 769.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER ME3 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER ME2 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER ME1 ;
  RECT 756.800 0.000 760.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER ME3 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER ME2 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER ME1 ;
  RECT 748.120 0.000 751.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER ME3 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER ME2 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER ME1 ;
  RECT 726.420 0.000 729.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 713.400 0.000 716.940 1.120 ;
  LAYER ME3 ;
  RECT 713.400 0.000 716.940 1.120 ;
  LAYER ME2 ;
  RECT 713.400 0.000 716.940 1.120 ;
  LAYER ME1 ;
  RECT 713.400 0.000 716.940 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER ME3 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER ME2 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER ME1 ;
  RECT 704.720 0.000 708.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER ME3 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER ME2 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER ME1 ;
  RECT 643.960 0.000 647.500 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER ME3 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER ME2 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER ME1 ;
  RECT 635.280 0.000 638.820 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER ME3 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER ME2 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER ME1 ;
  RECT 613.580 0.000 617.120 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER ME3 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER ME2 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER ME1 ;
  RECT 600.560 0.000 604.100 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER ME3 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER ME2 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER ME1 ;
  RECT 591.880 0.000 595.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER ME3 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER ME2 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER ME1 ;
  RECT 583.200 0.000 586.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER ME3 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER ME2 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER ME1 ;
  RECT 472.220 0.000 475.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER ME3 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER ME2 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER ME1 ;
  RECT 457.340 0.000 460.880 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER ME3 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER ME2 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER ME1 ;
  RECT 448.660 0.000 452.200 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER ME3 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER ME2 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER ME1 ;
  RECT 439.980 0.000 443.520 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER ME3 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER ME2 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER ME1 ;
  RECT 431.300 0.000 434.840 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.600 0.000 413.140 1.120 ;
  LAYER ME3 ;
  RECT 409.600 0.000 413.140 1.120 ;
  LAYER ME2 ;
  RECT 409.600 0.000 413.140 1.120 ;
  LAYER ME1 ;
  RECT 409.600 0.000 413.140 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.500 0.000 348.040 1.120 ;
  LAYER ME3 ;
  RECT 344.500 0.000 348.040 1.120 ;
  LAYER ME2 ;
  RECT 344.500 0.000 348.040 1.120 ;
  LAYER ME1 ;
  RECT 344.500 0.000 348.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.820 0.000 339.360 1.120 ;
  LAYER ME3 ;
  RECT 335.820 0.000 339.360 1.120 ;
  LAYER ME2 ;
  RECT 335.820 0.000 339.360 1.120 ;
  LAYER ME1 ;
  RECT 335.820 0.000 339.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.140 0.000 330.680 1.120 ;
  LAYER ME3 ;
  RECT 327.140 0.000 330.680 1.120 ;
  LAYER ME2 ;
  RECT 327.140 0.000 330.680 1.120 ;
  LAYER ME1 ;
  RECT 327.140 0.000 330.680 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME3 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME2 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME1 ;
  RECT 318.460 0.000 322.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME3 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME2 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME1 ;
  RECT 296.760 0.000 300.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER ME3 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER ME2 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER ME1 ;
  RECT 218.020 0.000 221.560 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.340 0.000 212.880 1.120 ;
  LAYER ME3 ;
  RECT 209.340 0.000 212.880 1.120 ;
  LAYER ME2 ;
  RECT 209.340 0.000 212.880 1.120 ;
  LAYER ME1 ;
  RECT 209.340 0.000 212.880 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.940 0.000 200.480 1.120 ;
  LAYER ME3 ;
  RECT 196.940 0.000 200.480 1.120 ;
  LAYER ME2 ;
  RECT 196.940 0.000 200.480 1.120 ;
  LAYER ME1 ;
  RECT 196.940 0.000 200.480 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER ME3 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER ME2 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER ME1 ;
  RECT 174.620 0.000 178.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER ME3 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER ME2 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER ME1 ;
  RECT 165.940 0.000 169.480 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER ME3 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER ME2 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER ME1 ;
  RECT 157.260 0.000 160.800 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.500 0.000 100.040 1.120 ;
  LAYER ME3 ;
  RECT 96.500 0.000 100.040 1.120 ;
  LAYER ME2 ;
  RECT 96.500 0.000 100.040 1.120 ;
  LAYER ME1 ;
  RECT 96.500 0.000 100.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER ME3 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER ME2 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER ME1 ;
  RECT 61.780 0.000 65.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER ME3 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER ME2 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER ME1 ;
  RECT 53.100 0.000 56.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER ME3 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER ME2 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER ME1 ;
  RECT 44.420 0.000 47.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
END GND
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 972.220 0.000 973.340 1.120 ;
  LAYER ME3 ;
  RECT 972.220 0.000 973.340 1.120 ;
  LAYER ME2 ;
  RECT 972.220 0.000 973.340 1.120 ;
  LAYER ME1 ;
  RECT 972.220 0.000 973.340 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 963.540 0.000 964.660 1.120 ;
  LAYER ME3 ;
  RECT 963.540 0.000 964.660 1.120 ;
  LAYER ME2 ;
  RECT 963.540 0.000 964.660 1.120 ;
  LAYER ME1 ;
  RECT 963.540 0.000 964.660 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 959.200 0.000 960.320 1.120 ;
  LAYER ME3 ;
  RECT 959.200 0.000 960.320 1.120 ;
  LAYER ME2 ;
  RECT 959.200 0.000 960.320 1.120 ;
  LAYER ME1 ;
  RECT 959.200 0.000 960.320 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 950.520 0.000 951.640 1.120 ;
  LAYER ME3 ;
  RECT 950.520 0.000 951.640 1.120 ;
  LAYER ME2 ;
  RECT 950.520 0.000 951.640 1.120 ;
  LAYER ME1 ;
  RECT 950.520 0.000 951.640 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 915.800 0.000 916.920 1.120 ;
  LAYER ME3 ;
  RECT 915.800 0.000 916.920 1.120 ;
  LAYER ME2 ;
  RECT 915.800 0.000 916.920 1.120 ;
  LAYER ME1 ;
  RECT 915.800 0.000 916.920 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 907.120 0.000 908.240 1.120 ;
  LAYER ME3 ;
  RECT 907.120 0.000 908.240 1.120 ;
  LAYER ME2 ;
  RECT 907.120 0.000 908.240 1.120 ;
  LAYER ME1 ;
  RECT 907.120 0.000 908.240 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 902.160 0.000 903.280 1.120 ;
  LAYER ME3 ;
  RECT 902.160 0.000 903.280 1.120 ;
  LAYER ME2 ;
  RECT 902.160 0.000 903.280 1.120 ;
  LAYER ME1 ;
  RECT 902.160 0.000 903.280 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 894.100 0.000 895.220 1.120 ;
  LAYER ME3 ;
  RECT 894.100 0.000 895.220 1.120 ;
  LAYER ME2 ;
  RECT 894.100 0.000 895.220 1.120 ;
  LAYER ME1 ;
  RECT 894.100 0.000 895.220 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME3 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME2 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME1 ;
  RECT 859.380 0.000 860.500 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 850.700 0.000 851.820 1.120 ;
  LAYER ME3 ;
  RECT 850.700 0.000 851.820 1.120 ;
  LAYER ME2 ;
  RECT 850.700 0.000 851.820 1.120 ;
  LAYER ME1 ;
  RECT 850.700 0.000 851.820 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER ME3 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER ME2 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER ME1 ;
  RECT 845.740 0.000 846.860 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 837.680 0.000 838.800 1.120 ;
  LAYER ME3 ;
  RECT 837.680 0.000 838.800 1.120 ;
  LAYER ME2 ;
  RECT 837.680 0.000 838.800 1.120 ;
  LAYER ME1 ;
  RECT 837.680 0.000 838.800 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER ME3 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER ME2 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER ME1 ;
  RECT 802.340 0.000 803.460 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 794.280 0.000 795.400 1.120 ;
  LAYER ME3 ;
  RECT 794.280 0.000 795.400 1.120 ;
  LAYER ME2 ;
  RECT 794.280 0.000 795.400 1.120 ;
  LAYER ME1 ;
  RECT 794.280 0.000 795.400 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 789.320 0.000 790.440 1.120 ;
  LAYER ME3 ;
  RECT 789.320 0.000 790.440 1.120 ;
  LAYER ME2 ;
  RECT 789.320 0.000 790.440 1.120 ;
  LAYER ME1 ;
  RECT 789.320 0.000 790.440 1.120 ;
 END
END DO24
PIN WEB3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 784.980 0.000 786.100 1.120 ;
  LAYER ME3 ;
  RECT 784.980 0.000 786.100 1.120 ;
  LAYER ME2 ;
  RECT 784.980 0.000 786.100 1.120 ;
  LAYER ME1 ;
  RECT 784.980 0.000 786.100 1.120 ;
 END
END WEB3
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER ME3 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER ME2 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER ME1 ;
  RECT 781.260 0.000 782.380 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 745.920 0.000 747.040 1.120 ;
  LAYER ME3 ;
  RECT 745.920 0.000 747.040 1.120 ;
  LAYER ME2 ;
  RECT 745.920 0.000 747.040 1.120 ;
  LAYER ME1 ;
  RECT 745.920 0.000 747.040 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 737.860 0.000 738.980 1.120 ;
  LAYER ME3 ;
  RECT 737.860 0.000 738.980 1.120 ;
  LAYER ME2 ;
  RECT 737.860 0.000 738.980 1.120 ;
  LAYER ME1 ;
  RECT 737.860 0.000 738.980 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME3 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME2 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME1 ;
  RECT 732.900 0.000 734.020 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 724.220 0.000 725.340 1.120 ;
  LAYER ME3 ;
  RECT 724.220 0.000 725.340 1.120 ;
  LAYER ME2 ;
  RECT 724.220 0.000 725.340 1.120 ;
  LAYER ME1 ;
  RECT 724.220 0.000 725.340 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 689.500 0.000 690.620 1.120 ;
  LAYER ME3 ;
  RECT 689.500 0.000 690.620 1.120 ;
  LAYER ME2 ;
  RECT 689.500 0.000 690.620 1.120 ;
  LAYER ME1 ;
  RECT 689.500 0.000 690.620 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 681.440 0.000 682.560 1.120 ;
  LAYER ME3 ;
  RECT 681.440 0.000 682.560 1.120 ;
  LAYER ME2 ;
  RECT 681.440 0.000 682.560 1.120 ;
  LAYER ME1 ;
  RECT 681.440 0.000 682.560 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME3 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME2 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME1 ;
  RECT 676.480 0.000 677.600 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 667.800 0.000 668.920 1.120 ;
  LAYER ME3 ;
  RECT 667.800 0.000 668.920 1.120 ;
  LAYER ME2 ;
  RECT 667.800 0.000 668.920 1.120 ;
  LAYER ME1 ;
  RECT 667.800 0.000 668.920 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 633.080 0.000 634.200 1.120 ;
  LAYER ME3 ;
  RECT 633.080 0.000 634.200 1.120 ;
  LAYER ME2 ;
  RECT 633.080 0.000 634.200 1.120 ;
  LAYER ME1 ;
  RECT 633.080 0.000 634.200 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 624.400 0.000 625.520 1.120 ;
  LAYER ME3 ;
  RECT 624.400 0.000 625.520 1.120 ;
  LAYER ME2 ;
  RECT 624.400 0.000 625.520 1.120 ;
  LAYER ME1 ;
  RECT 624.400 0.000 625.520 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME3 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME2 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME1 ;
  RECT 620.060 0.000 621.180 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 611.380 0.000 612.500 1.120 ;
  LAYER ME3 ;
  RECT 611.380 0.000 612.500 1.120 ;
  LAYER ME2 ;
  RECT 611.380 0.000 612.500 1.120 ;
  LAYER ME1 ;
  RECT 611.380 0.000 612.500 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME3 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME2 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME1 ;
  RECT 576.660 0.000 577.780 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 567.980 0.000 569.100 1.120 ;
  LAYER ME3 ;
  RECT 567.980 0.000 569.100 1.120 ;
  LAYER ME2 ;
  RECT 567.980 0.000 569.100 1.120 ;
  LAYER ME1 ;
  RECT 567.980 0.000 569.100 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 563.020 0.000 564.140 1.120 ;
  LAYER ME3 ;
  RECT 563.020 0.000 564.140 1.120 ;
  LAYER ME2 ;
  RECT 563.020 0.000 564.140 1.120 ;
  LAYER ME1 ;
  RECT 563.020 0.000 564.140 1.120 ;
 END
END DO16
PIN WEB2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 558.680 0.000 559.800 1.120 ;
  LAYER ME3 ;
  RECT 558.680 0.000 559.800 1.120 ;
  LAYER ME2 ;
  RECT 558.680 0.000 559.800 1.120 ;
  LAYER ME1 ;
  RECT 558.680 0.000 559.800 1.120 ;
 END
END WEB2
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 554.960 0.000 556.080 1.120 ;
  LAYER ME3 ;
  RECT 554.960 0.000 556.080 1.120 ;
  LAYER ME2 ;
  RECT 554.960 0.000 556.080 1.120 ;
  LAYER ME1 ;
  RECT 554.960 0.000 556.080 1.120 ;
 END
END DI16
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 548.760 0.000 549.880 1.120 ;
  LAYER ME3 ;
  RECT 548.760 0.000 549.880 1.120 ;
  LAYER ME2 ;
  RECT 548.760 0.000 549.880 1.120 ;
  LAYER ME1 ;
  RECT 548.760 0.000 549.880 1.120 ;
 END
END A1
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 542.560 0.000 543.680 1.120 ;
  LAYER ME3 ;
  RECT 542.560 0.000 543.680 1.120 ;
  LAYER ME2 ;
  RECT 542.560 0.000 543.680 1.120 ;
  LAYER ME1 ;
  RECT 542.560 0.000 543.680 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 540.700 0.000 541.820 1.120 ;
  LAYER ME3 ;
  RECT 540.700 0.000 541.820 1.120 ;
  LAYER ME2 ;
  RECT 540.700 0.000 541.820 1.120 ;
  LAYER ME1 ;
  RECT 540.700 0.000 541.820 1.120 ;
 END
END CS
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER ME3 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER ME2 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER ME1 ;
  RECT 538.840 0.000 539.960 1.120 ;
 END
END A3
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 519.000 0.000 520.120 1.120 ;
  LAYER ME3 ;
  RECT 519.000 0.000 520.120 1.120 ;
  LAYER ME2 ;
  RECT 519.000 0.000 520.120 1.120 ;
  LAYER ME1 ;
  RECT 519.000 0.000 520.120 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 515.900 0.000 517.020 1.120 ;
  LAYER ME3 ;
  RECT 515.900 0.000 517.020 1.120 ;
  LAYER ME2 ;
  RECT 515.900 0.000 517.020 1.120 ;
  LAYER ME1 ;
  RECT 515.900 0.000 517.020 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 514.040 0.000 515.160 1.120 ;
  LAYER ME3 ;
  RECT 514.040 0.000 515.160 1.120 ;
  LAYER ME2 ;
  RECT 514.040 0.000 515.160 1.120 ;
  LAYER ME1 ;
  RECT 514.040 0.000 515.160 1.120 ;
 END
END A0
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME3 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME2 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME1 ;
  RECT 509.700 0.000 510.820 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 501.640 0.000 502.760 1.120 ;
  LAYER ME3 ;
  RECT 501.640 0.000 502.760 1.120 ;
  LAYER ME2 ;
  RECT 501.640 0.000 502.760 1.120 ;
  LAYER ME1 ;
  RECT 501.640 0.000 502.760 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER ME3 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER ME2 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER ME1 ;
  RECT 499.160 0.000 500.280 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER ME3 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER ME2 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER ME1 ;
  RECT 491.100 0.000 492.220 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END A8
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER ME3 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER ME2 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER ME1 ;
  RECT 480.560 0.000 481.680 1.120 ;
 END
END A9
PIN A10
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME3 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME2 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME1 ;
  RECT 477.460 0.000 478.580 1.120 ;
 END
END A10
PIN A11
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER ME3 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER ME2 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER ME1 ;
  RECT 470.020 0.000 471.140 1.120 ;
 END
END A11
PIN A12
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 466.920 0.000 468.040 1.120 ;
  LAYER ME3 ;
  RECT 466.920 0.000 468.040 1.120 ;
  LAYER ME2 ;
  RECT 466.920 0.000 468.040 1.120 ;
  LAYER ME1 ;
  RECT 466.920 0.000 468.040 1.120 ;
 END
END A12
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME3 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME2 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME1 ;
  RECT 420.420 0.000 421.540 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME3 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME2 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME1 ;
  RECT 415.460 0.000 416.580 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME3 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME2 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME1 ;
  RECT 407.400 0.000 408.520 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME3 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME2 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME1 ;
  RECT 372.680 0.000 373.800 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME3 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME2 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME1 ;
  RECT 364.000 0.000 365.120 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME3 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME2 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME1 ;
  RECT 350.980 0.000 352.100 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME3 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME2 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME1 ;
  RECT 316.260 0.000 317.380 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME3 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME2 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME1 ;
  RECT 307.580 0.000 308.700 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME3 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME2 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME1 ;
  RECT 302.620 0.000 303.740 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME3 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME2 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME1 ;
  RECT 294.560 0.000 295.680 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO8
PIN WEB1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 241.860 0.000 242.980 1.120 ;
  LAYER ME3 ;
  RECT 241.860 0.000 242.980 1.120 ;
  LAYER ME2 ;
  RECT 241.860 0.000 242.980 1.120 ;
  LAYER ME1 ;
  RECT 241.860 0.000 242.980 1.120 ;
 END
END WEB1
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN WEB0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER ME3 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER ME2 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER ME1 ;
  RECT 15.560 0.000 16.680 1.120 ;
 END
END WEB0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 1015.560 1391.600 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 1015.560 1391.600 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 1015.560 1391.600 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 1015.560 1391.600 ;
  LAYER VI1 ;
  RECT 0.000 0.140 1015.560 1391.600 ;
  LAYER VI2 ;
  RECT 0.000 0.140 1015.560 1391.600 ;
  LAYER VI3 ;
  RECT 0.000 0.140 1015.560 1391.600 ;
END
END SUMA180_8192X8X4BM2
END LIBRARY



