parameter [1:0] ALU_SRC_RS        = 2'b00,
                ALU_SRC_EX_MEM_RD = 2'b01,
                ALU_SRC_MEM_WB_RD = 2'b10;

parameter       DATA_SRC_RS = 1'b0,
                DATA_SRC_RD = 1'b1;
