AHB/Decoder.sv