AHB/DefaultSlave.sv