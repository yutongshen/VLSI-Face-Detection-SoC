AHB/Arbiter.sv