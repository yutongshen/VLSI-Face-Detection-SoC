../include/def.svh