PLIC/Gateway.sv